VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_32x8
  FOREIGN sram_32x8 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 160.000 BY 2000.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.400 1.200 80.600 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.400 1.200 96.600 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.400 1.200 112.600 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.400 1.200 128.600 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.400 1.200 144.600 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 159.400 1.200 160.600 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.400 1.200 176.600 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 191.400 1.200 192.600 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 207.400 1.200 208.600 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.400 1.200 224.600 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 239.400 1.200 240.600 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 255.400 1.200 256.600 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 271.400 1.200 272.600 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 287.400 1.200 288.600 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 303.400 1.200 304.600 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 319.400 1.200 320.600 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 335.400 1.200 336.600 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 351.400 1.200 352.600 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 367.400 1.200 368.600 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 383.400 1.200 384.600 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.400 1.200 400.600 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 415.400 1.200 416.600 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 431.400 1.200 432.600 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 447.400 1.200 448.600 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 463.400 1.200 464.600 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 479.400 1.200 480.600 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 495.400 1.200 496.600 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 511.400 1.200 512.600 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 527.400 1.200 528.600 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.400 1.200 544.600 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 559.400 1.200 560.600 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 575.400 1.200 576.600 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 615.400 1.200 616.600 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 631.400 1.200 632.600 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 647.400 1.200 648.600 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 663.400 1.200 664.600 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 679.400 1.200 680.600 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 695.400 1.200 696.600 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 711.400 1.200 712.600 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 727.400 1.200 728.600 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 743.400 1.200 744.600 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 759.400 1.200 760.600 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 775.400 1.200 776.600 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 791.400 1.200 792.600 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 807.400 1.200 808.600 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 823.400 1.200 824.600 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 839.400 1.200 840.600 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 855.400 1.200 856.600 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 871.400 1.200 872.600 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 887.400 1.200 888.600 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 903.400 1.200 904.600 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 919.400 1.200 920.600 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 935.400 1.200 936.600 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 951.400 1.200 952.600 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 967.400 1.200 968.600 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 983.400 1.200 984.600 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 999.400 1.200 1000.600 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1015.400 1.200 1016.600 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1031.400 1.200 1032.600 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1047.400 1.200 1048.600 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1063.400 1.200 1064.600 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1079.400 1.200 1080.600 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1095.400 1.200 1096.600 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1111.400 1.200 1112.600 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1151.400 1.200 1152.600 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1167.400 1.200 1168.600 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1183.400 1.200 1184.600 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1199.400 1.200 1200.600 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1215.400 1.200 1216.600 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1231.400 1.200 1232.600 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1247.400 1.200 1248.600 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1263.400 1.200 1264.600 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1279.400 1.200 1280.600 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1295.400 1.200 1296.600 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1311.400 1.200 1312.600 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1327.400 1.200 1328.600 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1343.400 1.200 1344.600 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1359.400 1.200 1360.600 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1375.400 1.200 1376.600 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1391.400 1.200 1392.600 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1407.400 1.200 1408.600 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1423.400 1.200 1424.600 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1439.400 1.200 1440.600 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1455.400 1.200 1456.600 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1471.400 1.200 1472.600 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1487.400 1.200 1488.600 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1503.400 1.200 1504.600 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1519.400 1.200 1520.600 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1535.400 1.200 1536.600 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1551.400 1.200 1552.600 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1567.400 1.200 1568.600 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1583.400 1.200 1584.600 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1599.400 1.200 1600.600 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1615.400 1.200 1616.600 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1631.400 1.200 1632.600 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1647.400 1.200 1648.600 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1687.400 1.200 1688.600 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1703.400 1.200 1704.600 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1719.400 1.200 1720.600 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1735.400 1.200 1736.600 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1751.400 1.200 1752.600 ;
    END
  END addr_in[4]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1791.400 1.200 1792.600 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1807.400 1.200 1808.600 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 1823.400 1.200 1824.600 ;
    END
  END clk
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 77.600 80.000 82.400 1920.000 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
    END
  END vccd1
  OBS
    LAYER met1 ;
    RECT 0 0 160.000 2000.000 ;
    LAYER met2 ;
    RECT 0 0 160.000 2000.000 ;
    LAYER met3 ;
    RECT 1.200 0 160.000 2000.000 ;
    RECT 0 0.000 1.200 79.400 ;
    RECT 0 80.600 1.200 95.400 ;
    RECT 0 96.600 1.200 111.400 ;
    RECT 0 112.600 1.200 127.400 ;
    RECT 0 128.600 1.200 143.400 ;
    RECT 0 144.600 1.200 159.400 ;
    RECT 0 160.600 1.200 175.400 ;
    RECT 0 176.600 1.200 191.400 ;
    RECT 0 192.600 1.200 207.400 ;
    RECT 0 208.600 1.200 223.400 ;
    RECT 0 224.600 1.200 239.400 ;
    RECT 0 240.600 1.200 255.400 ;
    RECT 0 256.600 1.200 271.400 ;
    RECT 0 272.600 1.200 287.400 ;
    RECT 0 288.600 1.200 303.400 ;
    RECT 0 304.600 1.200 319.400 ;
    RECT 0 320.600 1.200 335.400 ;
    RECT 0 336.600 1.200 351.400 ;
    RECT 0 352.600 1.200 367.400 ;
    RECT 0 368.600 1.200 383.400 ;
    RECT 0 384.600 1.200 399.400 ;
    RECT 0 400.600 1.200 415.400 ;
    RECT 0 416.600 1.200 431.400 ;
    RECT 0 432.600 1.200 447.400 ;
    RECT 0 448.600 1.200 463.400 ;
    RECT 0 464.600 1.200 479.400 ;
    RECT 0 480.600 1.200 495.400 ;
    RECT 0 496.600 1.200 511.400 ;
    RECT 0 512.600 1.200 527.400 ;
    RECT 0 528.600 1.200 543.400 ;
    RECT 0 544.600 1.200 559.400 ;
    RECT 0 560.600 1.200 575.400 ;
    RECT 0 576.600 1.200 615.400 ;
    RECT 0 616.600 1.200 631.400 ;
    RECT 0 632.600 1.200 647.400 ;
    RECT 0 648.600 1.200 663.400 ;
    RECT 0 664.600 1.200 679.400 ;
    RECT 0 680.600 1.200 695.400 ;
    RECT 0 696.600 1.200 711.400 ;
    RECT 0 712.600 1.200 727.400 ;
    RECT 0 728.600 1.200 743.400 ;
    RECT 0 744.600 1.200 759.400 ;
    RECT 0 760.600 1.200 775.400 ;
    RECT 0 776.600 1.200 791.400 ;
    RECT 0 792.600 1.200 807.400 ;
    RECT 0 808.600 1.200 823.400 ;
    RECT 0 824.600 1.200 839.400 ;
    RECT 0 840.600 1.200 855.400 ;
    RECT 0 856.600 1.200 871.400 ;
    RECT 0 872.600 1.200 887.400 ;
    RECT 0 888.600 1.200 903.400 ;
    RECT 0 904.600 1.200 919.400 ;
    RECT 0 920.600 1.200 935.400 ;
    RECT 0 936.600 1.200 951.400 ;
    RECT 0 952.600 1.200 967.400 ;
    RECT 0 968.600 1.200 983.400 ;
    RECT 0 984.600 1.200 999.400 ;
    RECT 0 1000.600 1.200 1015.400 ;
    RECT 0 1016.600 1.200 1031.400 ;
    RECT 0 1032.600 1.200 1047.400 ;
    RECT 0 1048.600 1.200 1063.400 ;
    RECT 0 1064.600 1.200 1079.400 ;
    RECT 0 1080.600 1.200 1095.400 ;
    RECT 0 1096.600 1.200 1111.400 ;
    RECT 0 1112.600 1.200 1151.400 ;
    RECT 0 1152.600 1.200 1167.400 ;
    RECT 0 1168.600 1.200 1183.400 ;
    RECT 0 1184.600 1.200 1199.400 ;
    RECT 0 1200.600 1.200 1215.400 ;
    RECT 0 1216.600 1.200 1231.400 ;
    RECT 0 1232.600 1.200 1247.400 ;
    RECT 0 1248.600 1.200 1263.400 ;
    RECT 0 1264.600 1.200 1279.400 ;
    RECT 0 1280.600 1.200 1295.400 ;
    RECT 0 1296.600 1.200 1311.400 ;
    RECT 0 1312.600 1.200 1327.400 ;
    RECT 0 1328.600 1.200 1343.400 ;
    RECT 0 1344.600 1.200 1359.400 ;
    RECT 0 1360.600 1.200 1375.400 ;
    RECT 0 1376.600 1.200 1391.400 ;
    RECT 0 1392.600 1.200 1407.400 ;
    RECT 0 1408.600 1.200 1423.400 ;
    RECT 0 1424.600 1.200 1439.400 ;
    RECT 0 1440.600 1.200 1455.400 ;
    RECT 0 1456.600 1.200 1471.400 ;
    RECT 0 1472.600 1.200 1487.400 ;
    RECT 0 1488.600 1.200 1503.400 ;
    RECT 0 1504.600 1.200 1519.400 ;
    RECT 0 1520.600 1.200 1535.400 ;
    RECT 0 1536.600 1.200 1551.400 ;
    RECT 0 1552.600 1.200 1567.400 ;
    RECT 0 1568.600 1.200 1583.400 ;
    RECT 0 1584.600 1.200 1599.400 ;
    RECT 0 1600.600 1.200 1615.400 ;
    RECT 0 1616.600 1.200 1631.400 ;
    RECT 0 1632.600 1.200 1647.400 ;
    RECT 0 1648.600 1.200 1687.400 ;
    RECT 0 1688.600 1.200 1703.400 ;
    RECT 0 1704.600 1.200 1719.400 ;
    RECT 0 1720.600 1.200 1735.400 ;
    RECT 0 1736.600 1.200 1751.400 ;
    RECT 0 1752.600 1.200 1791.400 ;
    RECT 0 1792.600 1.200 1807.400 ;
    RECT 0 1808.600 1.200 1823.400 ;
    RECT 0 1824.600 1.200 2000.000 ;
    LAYER met4 ;
    RECT 0 0 160.000 80.000 ;
    RECT 0 1920.000 160.000 2000.000 ;
    RECT 0.000 80.000 77.600 1920.000 ;
    RECT 82.400 80.000 160.000 1920.000 ;
  END
END sram_32x8

END LIBRARY
