

module bsg_dff_width_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p7
(
  clk_i,
  data_i,
  data_o
);

  input [6:0] data_i;
  output [6:0] data_o;
  input clk_i;
  wire [6:0] data_o;
  reg data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_circular_ptr_slots_p3_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] o,n_o,ptr_nowrap;
  wire N0,N1,N2,N3,N4,N5;
  wire [2:0] ptr_wrap;
  reg o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign ptr_nowrap = o + add_i[0];
  assign { N4, N3, N2 } = o - { 1'b1, 1'b1 };
  assign ptr_wrap = { N4, N3, N2 } + add_i[0];
  assign n_o = (N0)? ptr_wrap[1:0] : 
               (N1)? ptr_nowrap : 1'b0;
  assign N0 = N5;
  assign N1 = ptr_wrap[2];
  assign N5 = ~ptr_wrap[2];

  always @(posedge clk) begin
    if(reset_i) begin
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_els_p3
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,N0,N1,N2,enq_r,deq_r,N3,equal_ptrs,sv2v_dc_1,sv2v_dc_2;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_slots_p3_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p3_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N3 = (N0)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = N1;
  assign N1 = enq_i | deq_i;
  assign N2 = ~N1;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N3) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p97_els_p3_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [96:0] w_data_i;
  input [1:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  wire [290:0] \nz.mem ;
  reg \nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,
  \nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,
  \nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,
  \nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,
  \nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,
  \nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,
  \nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,
  \nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,
  \nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,
  \nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,
  \nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,
  \nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,
  \nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,
  \nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,
  \nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,
  \nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,
  \nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,
  \nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,
  \nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,
  \nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,
  \nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,
  \nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,
  \nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,
  \nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,
  \nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,
  \nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,
  \nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,
  \nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,
  \nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,
  \nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,
  \nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,
  \nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,
  \nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,
  \nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,
  \nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,
  \nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,
  \nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,
  \nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,
  \nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,
  \nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,
  \nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,
  \nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,
  \nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,
  \nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,
  \nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,
  \nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,
  \nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,
  \nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,
  \nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,
  \nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,
  \nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,
  \nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,
  \nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,
  \nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,
  \nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,
  \nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,
  \nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,
  \nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,
  \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,
  \nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N11 = N4 & N5;
  assign N4 = ~r_addr_i[0];
  assign N5 = ~r_addr_i[1];
  assign { N18, N17, N16 } = (N6)? { N15, N14, N13 } : 
                             (N7)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = w_v_i;
  assign N7 = N12;
  assign r_data_o[96] = (N8)? \nz.mem [96] : 
                        (N9)? \nz.mem [193] : 
                        (N10)? \nz.mem [290] : 1'b0;
  assign N8 = N11;
  assign N9 = r_addr_i[0];
  assign N10 = r_addr_i[1];
  assign r_data_o[95] = (N8)? \nz.mem [95] : 
                        (N9)? \nz.mem [192] : 
                        (N10)? \nz.mem [289] : 1'b0;
  assign r_data_o[94] = (N8)? \nz.mem [94] : 
                        (N9)? \nz.mem [191] : 
                        (N10)? \nz.mem [288] : 1'b0;
  assign r_data_o[93] = (N8)? \nz.mem [93] : 
                        (N9)? \nz.mem [190] : 
                        (N10)? \nz.mem [287] : 1'b0;
  assign r_data_o[92] = (N8)? \nz.mem [92] : 
                        (N9)? \nz.mem [189] : 
                        (N10)? \nz.mem [286] : 1'b0;
  assign r_data_o[91] = (N8)? \nz.mem [91] : 
                        (N9)? \nz.mem [188] : 
                        (N10)? \nz.mem [285] : 1'b0;
  assign r_data_o[90] = (N8)? \nz.mem [90] : 
                        (N9)? \nz.mem [187] : 
                        (N10)? \nz.mem [284] : 1'b0;
  assign r_data_o[89] = (N8)? \nz.mem [89] : 
                        (N9)? \nz.mem [186] : 
                        (N10)? \nz.mem [283] : 1'b0;
  assign r_data_o[88] = (N8)? \nz.mem [88] : 
                        (N9)? \nz.mem [185] : 
                        (N10)? \nz.mem [282] : 1'b0;
  assign r_data_o[87] = (N8)? \nz.mem [87] : 
                        (N9)? \nz.mem [184] : 
                        (N10)? \nz.mem [281] : 1'b0;
  assign r_data_o[86] = (N8)? \nz.mem [86] : 
                        (N9)? \nz.mem [183] : 
                        (N10)? \nz.mem [280] : 1'b0;
  assign r_data_o[85] = (N8)? \nz.mem [85] : 
                        (N9)? \nz.mem [182] : 
                        (N10)? \nz.mem [279] : 1'b0;
  assign r_data_o[84] = (N8)? \nz.mem [84] : 
                        (N9)? \nz.mem [181] : 
                        (N10)? \nz.mem [278] : 1'b0;
  assign r_data_o[83] = (N8)? \nz.mem [83] : 
                        (N9)? \nz.mem [180] : 
                        (N10)? \nz.mem [277] : 1'b0;
  assign r_data_o[82] = (N8)? \nz.mem [82] : 
                        (N9)? \nz.mem [179] : 
                        (N10)? \nz.mem [276] : 1'b0;
  assign r_data_o[81] = (N8)? \nz.mem [81] : 
                        (N9)? \nz.mem [178] : 
                        (N10)? \nz.mem [275] : 1'b0;
  assign r_data_o[80] = (N8)? \nz.mem [80] : 
                        (N9)? \nz.mem [177] : 
                        (N10)? \nz.mem [274] : 1'b0;
  assign r_data_o[79] = (N8)? \nz.mem [79] : 
                        (N9)? \nz.mem [176] : 
                        (N10)? \nz.mem [273] : 1'b0;
  assign r_data_o[78] = (N8)? \nz.mem [78] : 
                        (N9)? \nz.mem [175] : 
                        (N10)? \nz.mem [272] : 1'b0;
  assign r_data_o[77] = (N8)? \nz.mem [77] : 
                        (N9)? \nz.mem [174] : 
                        (N10)? \nz.mem [271] : 1'b0;
  assign r_data_o[76] = (N8)? \nz.mem [76] : 
                        (N9)? \nz.mem [173] : 
                        (N10)? \nz.mem [270] : 1'b0;
  assign r_data_o[75] = (N8)? \nz.mem [75] : 
                        (N9)? \nz.mem [172] : 
                        (N10)? \nz.mem [269] : 1'b0;
  assign r_data_o[74] = (N8)? \nz.mem [74] : 
                        (N9)? \nz.mem [171] : 
                        (N10)? \nz.mem [268] : 1'b0;
  assign r_data_o[73] = (N8)? \nz.mem [73] : 
                        (N9)? \nz.mem [170] : 
                        (N10)? \nz.mem [267] : 1'b0;
  assign r_data_o[72] = (N8)? \nz.mem [72] : 
                        (N9)? \nz.mem [169] : 
                        (N10)? \nz.mem [266] : 1'b0;
  assign r_data_o[71] = (N8)? \nz.mem [71] : 
                        (N9)? \nz.mem [168] : 
                        (N10)? \nz.mem [265] : 1'b0;
  assign r_data_o[70] = (N8)? \nz.mem [70] : 
                        (N9)? \nz.mem [167] : 
                        (N10)? \nz.mem [264] : 1'b0;
  assign r_data_o[69] = (N8)? \nz.mem [69] : 
                        (N9)? \nz.mem [166] : 
                        (N10)? \nz.mem [263] : 1'b0;
  assign r_data_o[68] = (N8)? \nz.mem [68] : 
                        (N9)? \nz.mem [165] : 
                        (N10)? \nz.mem [262] : 1'b0;
  assign r_data_o[67] = (N8)? \nz.mem [67] : 
                        (N9)? \nz.mem [164] : 
                        (N10)? \nz.mem [261] : 1'b0;
  assign r_data_o[66] = (N8)? \nz.mem [66] : 
                        (N9)? \nz.mem [163] : 
                        (N10)? \nz.mem [260] : 1'b0;
  assign r_data_o[65] = (N8)? \nz.mem [65] : 
                        (N9)? \nz.mem [162] : 
                        (N10)? \nz.mem [259] : 1'b0;
  assign r_data_o[64] = (N8)? \nz.mem [64] : 
                        (N9)? \nz.mem [161] : 
                        (N10)? \nz.mem [258] : 1'b0;
  assign r_data_o[63] = (N8)? \nz.mem [63] : 
                        (N9)? \nz.mem [160] : 
                        (N10)? \nz.mem [257] : 1'b0;
  assign r_data_o[62] = (N8)? \nz.mem [62] : 
                        (N9)? \nz.mem [159] : 
                        (N10)? \nz.mem [256] : 1'b0;
  assign r_data_o[61] = (N8)? \nz.mem [61] : 
                        (N9)? \nz.mem [158] : 
                        (N10)? \nz.mem [255] : 1'b0;
  assign r_data_o[60] = (N8)? \nz.mem [60] : 
                        (N9)? \nz.mem [157] : 
                        (N10)? \nz.mem [254] : 1'b0;
  assign r_data_o[59] = (N8)? \nz.mem [59] : 
                        (N9)? \nz.mem [156] : 
                        (N10)? \nz.mem [253] : 1'b0;
  assign r_data_o[58] = (N8)? \nz.mem [58] : 
                        (N9)? \nz.mem [155] : 
                        (N10)? \nz.mem [252] : 1'b0;
  assign r_data_o[57] = (N8)? \nz.mem [57] : 
                        (N9)? \nz.mem [154] : 
                        (N10)? \nz.mem [251] : 1'b0;
  assign r_data_o[56] = (N8)? \nz.mem [56] : 
                        (N9)? \nz.mem [153] : 
                        (N10)? \nz.mem [250] : 1'b0;
  assign r_data_o[55] = (N8)? \nz.mem [55] : 
                        (N9)? \nz.mem [152] : 
                        (N10)? \nz.mem [249] : 1'b0;
  assign r_data_o[54] = (N8)? \nz.mem [54] : 
                        (N9)? \nz.mem [151] : 
                        (N10)? \nz.mem [248] : 1'b0;
  assign r_data_o[53] = (N8)? \nz.mem [53] : 
                        (N9)? \nz.mem [150] : 
                        (N10)? \nz.mem [247] : 1'b0;
  assign r_data_o[52] = (N8)? \nz.mem [52] : 
                        (N9)? \nz.mem [149] : 
                        (N10)? \nz.mem [246] : 1'b0;
  assign r_data_o[51] = (N8)? \nz.mem [51] : 
                        (N9)? \nz.mem [148] : 
                        (N10)? \nz.mem [245] : 1'b0;
  assign r_data_o[50] = (N8)? \nz.mem [50] : 
                        (N9)? \nz.mem [147] : 
                        (N10)? \nz.mem [244] : 1'b0;
  assign r_data_o[49] = (N8)? \nz.mem [49] : 
                        (N9)? \nz.mem [146] : 
                        (N10)? \nz.mem [243] : 1'b0;
  assign r_data_o[48] = (N8)? \nz.mem [48] : 
                        (N9)? \nz.mem [145] : 
                        (N10)? \nz.mem [242] : 1'b0;
  assign r_data_o[47] = (N8)? \nz.mem [47] : 
                        (N9)? \nz.mem [144] : 
                        (N10)? \nz.mem [241] : 1'b0;
  assign r_data_o[46] = (N8)? \nz.mem [46] : 
                        (N9)? \nz.mem [143] : 
                        (N10)? \nz.mem [240] : 1'b0;
  assign r_data_o[45] = (N8)? \nz.mem [45] : 
                        (N9)? \nz.mem [142] : 
                        (N10)? \nz.mem [239] : 1'b0;
  assign r_data_o[44] = (N8)? \nz.mem [44] : 
                        (N9)? \nz.mem [141] : 
                        (N10)? \nz.mem [238] : 1'b0;
  assign r_data_o[43] = (N8)? \nz.mem [43] : 
                        (N9)? \nz.mem [140] : 
                        (N10)? \nz.mem [237] : 1'b0;
  assign r_data_o[42] = (N8)? \nz.mem [42] : 
                        (N9)? \nz.mem [139] : 
                        (N10)? \nz.mem [236] : 1'b0;
  assign r_data_o[41] = (N8)? \nz.mem [41] : 
                        (N9)? \nz.mem [138] : 
                        (N10)? \nz.mem [235] : 1'b0;
  assign r_data_o[40] = (N8)? \nz.mem [40] : 
                        (N9)? \nz.mem [137] : 
                        (N10)? \nz.mem [234] : 1'b0;
  assign r_data_o[39] = (N8)? \nz.mem [39] : 
                        (N9)? \nz.mem [136] : 
                        (N10)? \nz.mem [233] : 1'b0;
  assign r_data_o[38] = (N8)? \nz.mem [38] : 
                        (N9)? \nz.mem [135] : 
                        (N10)? \nz.mem [232] : 1'b0;
  assign r_data_o[37] = (N8)? \nz.mem [37] : 
                        (N9)? \nz.mem [134] : 
                        (N10)? \nz.mem [231] : 1'b0;
  assign r_data_o[36] = (N8)? \nz.mem [36] : 
                        (N9)? \nz.mem [133] : 
                        (N10)? \nz.mem [230] : 1'b0;
  assign r_data_o[35] = (N8)? \nz.mem [35] : 
                        (N9)? \nz.mem [132] : 
                        (N10)? \nz.mem [229] : 1'b0;
  assign r_data_o[34] = (N8)? \nz.mem [34] : 
                        (N9)? \nz.mem [131] : 
                        (N10)? \nz.mem [228] : 1'b0;
  assign r_data_o[33] = (N8)? \nz.mem [33] : 
                        (N9)? \nz.mem [130] : 
                        (N10)? \nz.mem [227] : 1'b0;
  assign r_data_o[32] = (N8)? \nz.mem [32] : 
                        (N9)? \nz.mem [129] : 
                        (N10)? \nz.mem [226] : 1'b0;
  assign r_data_o[31] = (N8)? \nz.mem [31] : 
                        (N9)? \nz.mem [128] : 
                        (N10)? \nz.mem [225] : 1'b0;
  assign r_data_o[30] = (N8)? \nz.mem [30] : 
                        (N9)? \nz.mem [127] : 
                        (N10)? \nz.mem [224] : 1'b0;
  assign r_data_o[29] = (N8)? \nz.mem [29] : 
                        (N9)? \nz.mem [126] : 
                        (N10)? \nz.mem [223] : 1'b0;
  assign r_data_o[28] = (N8)? \nz.mem [28] : 
                        (N9)? \nz.mem [125] : 
                        (N10)? \nz.mem [222] : 1'b0;
  assign r_data_o[27] = (N8)? \nz.mem [27] : 
                        (N9)? \nz.mem [124] : 
                        (N10)? \nz.mem [221] : 1'b0;
  assign r_data_o[26] = (N8)? \nz.mem [26] : 
                        (N9)? \nz.mem [123] : 
                        (N10)? \nz.mem [220] : 1'b0;
  assign r_data_o[25] = (N8)? \nz.mem [25] : 
                        (N9)? \nz.mem [122] : 
                        (N10)? \nz.mem [219] : 1'b0;
  assign r_data_o[24] = (N8)? \nz.mem [24] : 
                        (N9)? \nz.mem [121] : 
                        (N10)? \nz.mem [218] : 1'b0;
  assign r_data_o[23] = (N8)? \nz.mem [23] : 
                        (N9)? \nz.mem [120] : 
                        (N10)? \nz.mem [217] : 1'b0;
  assign r_data_o[22] = (N8)? \nz.mem [22] : 
                        (N9)? \nz.mem [119] : 
                        (N10)? \nz.mem [216] : 1'b0;
  assign r_data_o[21] = (N8)? \nz.mem [21] : 
                        (N9)? \nz.mem [118] : 
                        (N10)? \nz.mem [215] : 1'b0;
  assign r_data_o[20] = (N8)? \nz.mem [20] : 
                        (N9)? \nz.mem [117] : 
                        (N10)? \nz.mem [214] : 1'b0;
  assign r_data_o[19] = (N8)? \nz.mem [19] : 
                        (N9)? \nz.mem [116] : 
                        (N10)? \nz.mem [213] : 1'b0;
  assign r_data_o[18] = (N8)? \nz.mem [18] : 
                        (N9)? \nz.mem [115] : 
                        (N10)? \nz.mem [212] : 1'b0;
  assign r_data_o[17] = (N8)? \nz.mem [17] : 
                        (N9)? \nz.mem [114] : 
                        (N10)? \nz.mem [211] : 1'b0;
  assign r_data_o[16] = (N8)? \nz.mem [16] : 
                        (N9)? \nz.mem [113] : 
                        (N10)? \nz.mem [210] : 1'b0;
  assign r_data_o[15] = (N8)? \nz.mem [15] : 
                        (N9)? \nz.mem [112] : 
                        (N10)? \nz.mem [209] : 1'b0;
  assign r_data_o[14] = (N8)? \nz.mem [14] : 
                        (N9)? \nz.mem [111] : 
                        (N10)? \nz.mem [208] : 1'b0;
  assign r_data_o[13] = (N8)? \nz.mem [13] : 
                        (N9)? \nz.mem [110] : 
                        (N10)? \nz.mem [207] : 1'b0;
  assign r_data_o[12] = (N8)? \nz.mem [12] : 
                        (N9)? \nz.mem [109] : 
                        (N10)? \nz.mem [206] : 1'b0;
  assign r_data_o[11] = (N8)? \nz.mem [11] : 
                        (N9)? \nz.mem [108] : 
                        (N10)? \nz.mem [205] : 1'b0;
  assign r_data_o[10] = (N8)? \nz.mem [10] : 
                        (N9)? \nz.mem [107] : 
                        (N10)? \nz.mem [204] : 1'b0;
  assign r_data_o[9] = (N8)? \nz.mem [9] : 
                       (N9)? \nz.mem [106] : 
                       (N10)? \nz.mem [203] : 1'b0;
  assign r_data_o[8] = (N8)? \nz.mem [8] : 
                       (N9)? \nz.mem [105] : 
                       (N10)? \nz.mem [202] : 1'b0;
  assign r_data_o[7] = (N8)? \nz.mem [7] : 
                       (N9)? \nz.mem [104] : 
                       (N10)? \nz.mem [201] : 1'b0;
  assign r_data_o[6] = (N8)? \nz.mem [6] : 
                       (N9)? \nz.mem [103] : 
                       (N10)? \nz.mem [200] : 1'b0;
  assign r_data_o[5] = (N8)? \nz.mem [5] : 
                       (N9)? \nz.mem [102] : 
                       (N10)? \nz.mem [199] : 1'b0;
  assign r_data_o[4] = (N8)? \nz.mem [4] : 
                       (N9)? \nz.mem [101] : 
                       (N10)? \nz.mem [198] : 1'b0;
  assign r_data_o[3] = (N8)? \nz.mem [3] : 
                       (N9)? \nz.mem [100] : 
                       (N10)? \nz.mem [197] : 1'b0;
  assign r_data_o[2] = (N8)? \nz.mem [2] : 
                       (N9)? \nz.mem [99] : 
                       (N10)? \nz.mem [196] : 1'b0;
  assign r_data_o[1] = (N8)? \nz.mem [1] : 
                       (N9)? \nz.mem [98] : 
                       (N10)? \nz.mem [195] : 1'b0;
  assign r_data_o[0] = (N8)? \nz.mem [0] : 
                       (N9)? \nz.mem [97] : 
                       (N10)? \nz.mem [194] : 1'b0;
  assign N12 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N18) begin
      \nz.mem_290_sv2v_reg  <= w_data_i[96];
      \nz.mem_289_sv2v_reg  <= w_data_i[95];
      \nz.mem_288_sv2v_reg  <= w_data_i[94];
      \nz.mem_287_sv2v_reg  <= w_data_i[93];
      \nz.mem_286_sv2v_reg  <= w_data_i[92];
      \nz.mem_285_sv2v_reg  <= w_data_i[91];
      \nz.mem_284_sv2v_reg  <= w_data_i[90];
      \nz.mem_283_sv2v_reg  <= w_data_i[89];
      \nz.mem_282_sv2v_reg  <= w_data_i[88];
      \nz.mem_281_sv2v_reg  <= w_data_i[87];
      \nz.mem_280_sv2v_reg  <= w_data_i[86];
      \nz.mem_279_sv2v_reg  <= w_data_i[85];
      \nz.mem_278_sv2v_reg  <= w_data_i[84];
      \nz.mem_277_sv2v_reg  <= w_data_i[83];
      \nz.mem_276_sv2v_reg  <= w_data_i[82];
      \nz.mem_275_sv2v_reg  <= w_data_i[81];
      \nz.mem_274_sv2v_reg  <= w_data_i[80];
      \nz.mem_273_sv2v_reg  <= w_data_i[79];
      \nz.mem_272_sv2v_reg  <= w_data_i[78];
      \nz.mem_271_sv2v_reg  <= w_data_i[77];
      \nz.mem_270_sv2v_reg  <= w_data_i[76];
      \nz.mem_269_sv2v_reg  <= w_data_i[75];
      \nz.mem_268_sv2v_reg  <= w_data_i[74];
      \nz.mem_267_sv2v_reg  <= w_data_i[73];
      \nz.mem_266_sv2v_reg  <= w_data_i[72];
      \nz.mem_265_sv2v_reg  <= w_data_i[71];
      \nz.mem_264_sv2v_reg  <= w_data_i[70];
      \nz.mem_263_sv2v_reg  <= w_data_i[69];
      \nz.mem_262_sv2v_reg  <= w_data_i[68];
      \nz.mem_261_sv2v_reg  <= w_data_i[67];
      \nz.mem_260_sv2v_reg  <= w_data_i[66];
      \nz.mem_259_sv2v_reg  <= w_data_i[65];
      \nz.mem_258_sv2v_reg  <= w_data_i[64];
      \nz.mem_257_sv2v_reg  <= w_data_i[63];
      \nz.mem_256_sv2v_reg  <= w_data_i[62];
      \nz.mem_255_sv2v_reg  <= w_data_i[61];
      \nz.mem_254_sv2v_reg  <= w_data_i[60];
      \nz.mem_253_sv2v_reg  <= w_data_i[59];
      \nz.mem_252_sv2v_reg  <= w_data_i[58];
      \nz.mem_251_sv2v_reg  <= w_data_i[57];
      \nz.mem_250_sv2v_reg  <= w_data_i[56];
      \nz.mem_249_sv2v_reg  <= w_data_i[55];
      \nz.mem_248_sv2v_reg  <= w_data_i[54];
      \nz.mem_247_sv2v_reg  <= w_data_i[53];
      \nz.mem_246_sv2v_reg  <= w_data_i[52];
      \nz.mem_245_sv2v_reg  <= w_data_i[51];
      \nz.mem_244_sv2v_reg  <= w_data_i[50];
      \nz.mem_243_sv2v_reg  <= w_data_i[49];
      \nz.mem_242_sv2v_reg  <= w_data_i[48];
      \nz.mem_241_sv2v_reg  <= w_data_i[47];
      \nz.mem_240_sv2v_reg  <= w_data_i[46];
      \nz.mem_239_sv2v_reg  <= w_data_i[45];
      \nz.mem_238_sv2v_reg  <= w_data_i[44];
      \nz.mem_237_sv2v_reg  <= w_data_i[43];
      \nz.mem_236_sv2v_reg  <= w_data_i[42];
      \nz.mem_235_sv2v_reg  <= w_data_i[41];
      \nz.mem_234_sv2v_reg  <= w_data_i[40];
      \nz.mem_233_sv2v_reg  <= w_data_i[39];
      \nz.mem_232_sv2v_reg  <= w_data_i[38];
      \nz.mem_231_sv2v_reg  <= w_data_i[37];
      \nz.mem_230_sv2v_reg  <= w_data_i[36];
      \nz.mem_229_sv2v_reg  <= w_data_i[35];
      \nz.mem_228_sv2v_reg  <= w_data_i[34];
      \nz.mem_227_sv2v_reg  <= w_data_i[33];
      \nz.mem_226_sv2v_reg  <= w_data_i[32];
      \nz.mem_225_sv2v_reg  <= w_data_i[31];
      \nz.mem_224_sv2v_reg  <= w_data_i[30];
      \nz.mem_223_sv2v_reg  <= w_data_i[29];
      \nz.mem_222_sv2v_reg  <= w_data_i[28];
      \nz.mem_221_sv2v_reg  <= w_data_i[27];
      \nz.mem_220_sv2v_reg  <= w_data_i[26];
      \nz.mem_219_sv2v_reg  <= w_data_i[25];
      \nz.mem_218_sv2v_reg  <= w_data_i[24];
      \nz.mem_217_sv2v_reg  <= w_data_i[23];
      \nz.mem_216_sv2v_reg  <= w_data_i[22];
      \nz.mem_215_sv2v_reg  <= w_data_i[21];
      \nz.mem_214_sv2v_reg  <= w_data_i[20];
      \nz.mem_213_sv2v_reg  <= w_data_i[19];
      \nz.mem_212_sv2v_reg  <= w_data_i[18];
      \nz.mem_211_sv2v_reg  <= w_data_i[17];
      \nz.mem_210_sv2v_reg  <= w_data_i[16];
      \nz.mem_209_sv2v_reg  <= w_data_i[15];
      \nz.mem_208_sv2v_reg  <= w_data_i[14];
      \nz.mem_207_sv2v_reg  <= w_data_i[13];
      \nz.mem_206_sv2v_reg  <= w_data_i[12];
      \nz.mem_205_sv2v_reg  <= w_data_i[11];
      \nz.mem_204_sv2v_reg  <= w_data_i[10];
      \nz.mem_203_sv2v_reg  <= w_data_i[9];
      \nz.mem_202_sv2v_reg  <= w_data_i[8];
      \nz.mem_201_sv2v_reg  <= w_data_i[7];
      \nz.mem_200_sv2v_reg  <= w_data_i[6];
      \nz.mem_199_sv2v_reg  <= w_data_i[5];
      \nz.mem_198_sv2v_reg  <= w_data_i[4];
      \nz.mem_197_sv2v_reg  <= w_data_i[3];
      \nz.mem_196_sv2v_reg  <= w_data_i[2];
      \nz.mem_195_sv2v_reg  <= w_data_i[1];
      \nz.mem_194_sv2v_reg  <= w_data_i[0];
    end 
    if(N17) begin
      \nz.mem_193_sv2v_reg  <= w_data_i[96];
      \nz.mem_192_sv2v_reg  <= w_data_i[95];
      \nz.mem_191_sv2v_reg  <= w_data_i[94];
      \nz.mem_190_sv2v_reg  <= w_data_i[93];
      \nz.mem_189_sv2v_reg  <= w_data_i[92];
      \nz.mem_188_sv2v_reg  <= w_data_i[91];
      \nz.mem_187_sv2v_reg  <= w_data_i[90];
      \nz.mem_186_sv2v_reg  <= w_data_i[89];
      \nz.mem_185_sv2v_reg  <= w_data_i[88];
      \nz.mem_184_sv2v_reg  <= w_data_i[87];
      \nz.mem_183_sv2v_reg  <= w_data_i[86];
      \nz.mem_182_sv2v_reg  <= w_data_i[85];
      \nz.mem_181_sv2v_reg  <= w_data_i[84];
      \nz.mem_180_sv2v_reg  <= w_data_i[83];
      \nz.mem_179_sv2v_reg  <= w_data_i[82];
      \nz.mem_178_sv2v_reg  <= w_data_i[81];
      \nz.mem_177_sv2v_reg  <= w_data_i[80];
      \nz.mem_176_sv2v_reg  <= w_data_i[79];
      \nz.mem_175_sv2v_reg  <= w_data_i[78];
      \nz.mem_174_sv2v_reg  <= w_data_i[77];
      \nz.mem_173_sv2v_reg  <= w_data_i[76];
      \nz.mem_172_sv2v_reg  <= w_data_i[75];
      \nz.mem_171_sv2v_reg  <= w_data_i[74];
      \nz.mem_170_sv2v_reg  <= w_data_i[73];
      \nz.mem_169_sv2v_reg  <= w_data_i[72];
      \nz.mem_168_sv2v_reg  <= w_data_i[71];
      \nz.mem_167_sv2v_reg  <= w_data_i[70];
      \nz.mem_166_sv2v_reg  <= w_data_i[69];
      \nz.mem_165_sv2v_reg  <= w_data_i[68];
      \nz.mem_164_sv2v_reg  <= w_data_i[67];
      \nz.mem_163_sv2v_reg  <= w_data_i[66];
      \nz.mem_162_sv2v_reg  <= w_data_i[65];
      \nz.mem_161_sv2v_reg  <= w_data_i[64];
      \nz.mem_160_sv2v_reg  <= w_data_i[63];
      \nz.mem_159_sv2v_reg  <= w_data_i[62];
      \nz.mem_158_sv2v_reg  <= w_data_i[61];
      \nz.mem_157_sv2v_reg  <= w_data_i[60];
      \nz.mem_156_sv2v_reg  <= w_data_i[59];
      \nz.mem_155_sv2v_reg  <= w_data_i[58];
      \nz.mem_154_sv2v_reg  <= w_data_i[57];
      \nz.mem_153_sv2v_reg  <= w_data_i[56];
      \nz.mem_152_sv2v_reg  <= w_data_i[55];
      \nz.mem_151_sv2v_reg  <= w_data_i[54];
      \nz.mem_150_sv2v_reg  <= w_data_i[53];
      \nz.mem_149_sv2v_reg  <= w_data_i[52];
      \nz.mem_148_sv2v_reg  <= w_data_i[51];
      \nz.mem_147_sv2v_reg  <= w_data_i[50];
      \nz.mem_146_sv2v_reg  <= w_data_i[49];
      \nz.mem_145_sv2v_reg  <= w_data_i[48];
      \nz.mem_144_sv2v_reg  <= w_data_i[47];
      \nz.mem_143_sv2v_reg  <= w_data_i[46];
      \nz.mem_142_sv2v_reg  <= w_data_i[45];
      \nz.mem_141_sv2v_reg  <= w_data_i[44];
      \nz.mem_140_sv2v_reg  <= w_data_i[43];
      \nz.mem_139_sv2v_reg  <= w_data_i[42];
      \nz.mem_138_sv2v_reg  <= w_data_i[41];
      \nz.mem_137_sv2v_reg  <= w_data_i[40];
      \nz.mem_136_sv2v_reg  <= w_data_i[39];
      \nz.mem_135_sv2v_reg  <= w_data_i[38];
      \nz.mem_134_sv2v_reg  <= w_data_i[37];
      \nz.mem_133_sv2v_reg  <= w_data_i[36];
      \nz.mem_132_sv2v_reg  <= w_data_i[35];
      \nz.mem_131_sv2v_reg  <= w_data_i[34];
      \nz.mem_130_sv2v_reg  <= w_data_i[33];
      \nz.mem_129_sv2v_reg  <= w_data_i[32];
      \nz.mem_128_sv2v_reg  <= w_data_i[31];
      \nz.mem_127_sv2v_reg  <= w_data_i[30];
      \nz.mem_126_sv2v_reg  <= w_data_i[29];
      \nz.mem_125_sv2v_reg  <= w_data_i[28];
      \nz.mem_124_sv2v_reg  <= w_data_i[27];
      \nz.mem_123_sv2v_reg  <= w_data_i[26];
      \nz.mem_122_sv2v_reg  <= w_data_i[25];
      \nz.mem_121_sv2v_reg  <= w_data_i[24];
      \nz.mem_120_sv2v_reg  <= w_data_i[23];
      \nz.mem_119_sv2v_reg  <= w_data_i[22];
      \nz.mem_118_sv2v_reg  <= w_data_i[21];
      \nz.mem_117_sv2v_reg  <= w_data_i[20];
      \nz.mem_116_sv2v_reg  <= w_data_i[19];
      \nz.mem_115_sv2v_reg  <= w_data_i[18];
      \nz.mem_114_sv2v_reg  <= w_data_i[17];
      \nz.mem_113_sv2v_reg  <= w_data_i[16];
      \nz.mem_112_sv2v_reg  <= w_data_i[15];
      \nz.mem_111_sv2v_reg  <= w_data_i[14];
      \nz.mem_110_sv2v_reg  <= w_data_i[13];
      \nz.mem_109_sv2v_reg  <= w_data_i[12];
      \nz.mem_108_sv2v_reg  <= w_data_i[11];
      \nz.mem_107_sv2v_reg  <= w_data_i[10];
      \nz.mem_106_sv2v_reg  <= w_data_i[9];
      \nz.mem_105_sv2v_reg  <= w_data_i[8];
      \nz.mem_104_sv2v_reg  <= w_data_i[7];
      \nz.mem_103_sv2v_reg  <= w_data_i[6];
      \nz.mem_102_sv2v_reg  <= w_data_i[5];
      \nz.mem_101_sv2v_reg  <= w_data_i[4];
      \nz.mem_100_sv2v_reg  <= w_data_i[3];
      \nz.mem_99_sv2v_reg  <= w_data_i[2];
      \nz.mem_98_sv2v_reg  <= w_data_i[1];
      \nz.mem_97_sv2v_reg  <= w_data_i[0];
    end 
    if(N16) begin
      \nz.mem_96_sv2v_reg  <= w_data_i[96];
      \nz.mem_95_sv2v_reg  <= w_data_i[95];
      \nz.mem_94_sv2v_reg  <= w_data_i[94];
      \nz.mem_93_sv2v_reg  <= w_data_i[93];
      \nz.mem_92_sv2v_reg  <= w_data_i[92];
      \nz.mem_91_sv2v_reg  <= w_data_i[91];
      \nz.mem_90_sv2v_reg  <= w_data_i[90];
      \nz.mem_89_sv2v_reg  <= w_data_i[89];
      \nz.mem_88_sv2v_reg  <= w_data_i[88];
      \nz.mem_87_sv2v_reg  <= w_data_i[87];
      \nz.mem_86_sv2v_reg  <= w_data_i[86];
      \nz.mem_85_sv2v_reg  <= w_data_i[85];
      \nz.mem_84_sv2v_reg  <= w_data_i[84];
      \nz.mem_83_sv2v_reg  <= w_data_i[83];
      \nz.mem_82_sv2v_reg  <= w_data_i[82];
      \nz.mem_81_sv2v_reg  <= w_data_i[81];
      \nz.mem_80_sv2v_reg  <= w_data_i[80];
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p97_els_p3_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [96:0] w_data_i;
  input [1:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;

  bsg_mem_1r1w_synth_width_p97_els_p3_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p97_els_p3_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [96:0] data_i;
  output [96:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [96:0] data_o;
  wire ready_o,v_o,enque,full,empty,sv2v_dc_1,sv2v_dc_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p3
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p97_els_p3_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_o;
  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p97_els_p3
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [96:0] data_i;
  output [96:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [96:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p97_els_p3_ready_THEN_valid_p0
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_dff_reset_width_p1_reset_val_p0
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p97_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [96:0] w_data_i;
  input [0:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [193:0] \nz.mem ;
  reg \nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,
  \nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,
  \nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,
  \nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,
  \nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,
  \nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,
  \nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,
  \nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,
  \nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,
  \nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,
  \nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,
  \nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,
  \nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,
  \nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,
  \nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,
  \nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,
  \nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,
  \nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,
  \nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,
  \nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,
  \nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,
  \nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,
  \nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,
  \nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,
  \nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,
  \nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,
  \nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,
  \nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,
  \nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,
  \nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,
  \nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,
  \nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,
  \nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,
  \nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,
  \nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,
  \nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,
  \nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,
  \nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,
  \nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,
  \nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[96] = (N3)? \nz.mem [96] : 
                        (N0)? \nz.mem [193] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[95] = (N3)? \nz.mem [95] : 
                        (N0)? \nz.mem [192] : 1'b0;
  assign r_data_o[94] = (N3)? \nz.mem [94] : 
                        (N0)? \nz.mem [191] : 1'b0;
  assign r_data_o[93] = (N3)? \nz.mem [93] : 
                        (N0)? \nz.mem [190] : 1'b0;
  assign r_data_o[92] = (N3)? \nz.mem [92] : 
                        (N0)? \nz.mem [189] : 1'b0;
  assign r_data_o[91] = (N3)? \nz.mem [91] : 
                        (N0)? \nz.mem [188] : 1'b0;
  assign r_data_o[90] = (N3)? \nz.mem [90] : 
                        (N0)? \nz.mem [187] : 1'b0;
  assign r_data_o[89] = (N3)? \nz.mem [89] : 
                        (N0)? \nz.mem [186] : 1'b0;
  assign r_data_o[88] = (N3)? \nz.mem [88] : 
                        (N0)? \nz.mem [185] : 1'b0;
  assign r_data_o[87] = (N3)? \nz.mem [87] : 
                        (N0)? \nz.mem [184] : 1'b0;
  assign r_data_o[86] = (N3)? \nz.mem [86] : 
                        (N0)? \nz.mem [183] : 1'b0;
  assign r_data_o[85] = (N3)? \nz.mem [85] : 
                        (N0)? \nz.mem [182] : 1'b0;
  assign r_data_o[84] = (N3)? \nz.mem [84] : 
                        (N0)? \nz.mem [181] : 1'b0;
  assign r_data_o[83] = (N3)? \nz.mem [83] : 
                        (N0)? \nz.mem [180] : 1'b0;
  assign r_data_o[82] = (N3)? \nz.mem [82] : 
                        (N0)? \nz.mem [179] : 1'b0;
  assign r_data_o[81] = (N3)? \nz.mem [81] : 
                        (N0)? \nz.mem [178] : 1'b0;
  assign r_data_o[80] = (N3)? \nz.mem [80] : 
                        (N0)? \nz.mem [177] : 1'b0;
  assign r_data_o[79] = (N3)? \nz.mem [79] : 
                        (N0)? \nz.mem [176] : 1'b0;
  assign r_data_o[78] = (N3)? \nz.mem [78] : 
                        (N0)? \nz.mem [175] : 1'b0;
  assign r_data_o[77] = (N3)? \nz.mem [77] : 
                        (N0)? \nz.mem [174] : 1'b0;
  assign r_data_o[76] = (N3)? \nz.mem [76] : 
                        (N0)? \nz.mem [173] : 1'b0;
  assign r_data_o[75] = (N3)? \nz.mem [75] : 
                        (N0)? \nz.mem [172] : 1'b0;
  assign r_data_o[74] = (N3)? \nz.mem [74] : 
                        (N0)? \nz.mem [171] : 1'b0;
  assign r_data_o[73] = (N3)? \nz.mem [73] : 
                        (N0)? \nz.mem [170] : 1'b0;
  assign r_data_o[72] = (N3)? \nz.mem [72] : 
                        (N0)? \nz.mem [169] : 1'b0;
  assign r_data_o[71] = (N3)? \nz.mem [71] : 
                        (N0)? \nz.mem [168] : 1'b0;
  assign r_data_o[70] = (N3)? \nz.mem [70] : 
                        (N0)? \nz.mem [167] : 1'b0;
  assign r_data_o[69] = (N3)? \nz.mem [69] : 
                        (N0)? \nz.mem [166] : 1'b0;
  assign r_data_o[68] = (N3)? \nz.mem [68] : 
                        (N0)? \nz.mem [165] : 1'b0;
  assign r_data_o[67] = (N3)? \nz.mem [67] : 
                        (N0)? \nz.mem [164] : 1'b0;
  assign r_data_o[66] = (N3)? \nz.mem [66] : 
                        (N0)? \nz.mem [163] : 1'b0;
  assign r_data_o[65] = (N3)? \nz.mem [65] : 
                        (N0)? \nz.mem [162] : 1'b0;
  assign r_data_o[64] = (N3)? \nz.mem [64] : 
                        (N0)? \nz.mem [161] : 1'b0;
  assign r_data_o[63] = (N3)? \nz.mem [63] : 
                        (N0)? \nz.mem [160] : 1'b0;
  assign r_data_o[62] = (N3)? \nz.mem [62] : 
                        (N0)? \nz.mem [159] : 1'b0;
  assign r_data_o[61] = (N3)? \nz.mem [61] : 
                        (N0)? \nz.mem [158] : 1'b0;
  assign r_data_o[60] = (N3)? \nz.mem [60] : 
                        (N0)? \nz.mem [157] : 1'b0;
  assign r_data_o[59] = (N3)? \nz.mem [59] : 
                        (N0)? \nz.mem [156] : 1'b0;
  assign r_data_o[58] = (N3)? \nz.mem [58] : 
                        (N0)? \nz.mem [155] : 1'b0;
  assign r_data_o[57] = (N3)? \nz.mem [57] : 
                        (N0)? \nz.mem [154] : 1'b0;
  assign r_data_o[56] = (N3)? \nz.mem [56] : 
                        (N0)? \nz.mem [153] : 1'b0;
  assign r_data_o[55] = (N3)? \nz.mem [55] : 
                        (N0)? \nz.mem [152] : 1'b0;
  assign r_data_o[54] = (N3)? \nz.mem [54] : 
                        (N0)? \nz.mem [151] : 1'b0;
  assign r_data_o[53] = (N3)? \nz.mem [53] : 
                        (N0)? \nz.mem [150] : 1'b0;
  assign r_data_o[52] = (N3)? \nz.mem [52] : 
                        (N0)? \nz.mem [149] : 1'b0;
  assign r_data_o[51] = (N3)? \nz.mem [51] : 
                        (N0)? \nz.mem [148] : 1'b0;
  assign r_data_o[50] = (N3)? \nz.mem [50] : 
                        (N0)? \nz.mem [147] : 1'b0;
  assign r_data_o[49] = (N3)? \nz.mem [49] : 
                        (N0)? \nz.mem [146] : 1'b0;
  assign r_data_o[48] = (N3)? \nz.mem [48] : 
                        (N0)? \nz.mem [145] : 1'b0;
  assign r_data_o[47] = (N3)? \nz.mem [47] : 
                        (N0)? \nz.mem [144] : 1'b0;
  assign r_data_o[46] = (N3)? \nz.mem [46] : 
                        (N0)? \nz.mem [143] : 1'b0;
  assign r_data_o[45] = (N3)? \nz.mem [45] : 
                        (N0)? \nz.mem [142] : 1'b0;
  assign r_data_o[44] = (N3)? \nz.mem [44] : 
                        (N0)? \nz.mem [141] : 1'b0;
  assign r_data_o[43] = (N3)? \nz.mem [43] : 
                        (N0)? \nz.mem [140] : 1'b0;
  assign r_data_o[42] = (N3)? \nz.mem [42] : 
                        (N0)? \nz.mem [139] : 1'b0;
  assign r_data_o[41] = (N3)? \nz.mem [41] : 
                        (N0)? \nz.mem [138] : 1'b0;
  assign r_data_o[40] = (N3)? \nz.mem [40] : 
                        (N0)? \nz.mem [137] : 1'b0;
  assign r_data_o[39] = (N3)? \nz.mem [39] : 
                        (N0)? \nz.mem [136] : 1'b0;
  assign r_data_o[38] = (N3)? \nz.mem [38] : 
                        (N0)? \nz.mem [135] : 1'b0;
  assign r_data_o[37] = (N3)? \nz.mem [37] : 
                        (N0)? \nz.mem [134] : 1'b0;
  assign r_data_o[36] = (N3)? \nz.mem [36] : 
                        (N0)? \nz.mem [133] : 1'b0;
  assign r_data_o[35] = (N3)? \nz.mem [35] : 
                        (N0)? \nz.mem [132] : 1'b0;
  assign r_data_o[34] = (N3)? \nz.mem [34] : 
                        (N0)? \nz.mem [131] : 1'b0;
  assign r_data_o[33] = (N3)? \nz.mem [33] : 
                        (N0)? \nz.mem [130] : 1'b0;
  assign r_data_o[32] = (N3)? \nz.mem [32] : 
                        (N0)? \nz.mem [129] : 1'b0;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [128] : 1'b0;
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [127] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [126] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [125] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [124] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [123] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [122] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [121] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [120] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [119] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [118] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [117] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [116] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [115] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [114] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [113] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [112] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [111] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [110] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [109] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [108] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [107] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [106] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [105] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [104] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [103] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [102] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [101] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [100] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [99] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [98] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [97] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_193_sv2v_reg  <= w_data_i[96];
      \nz.mem_192_sv2v_reg  <= w_data_i[95];
      \nz.mem_191_sv2v_reg  <= w_data_i[94];
      \nz.mem_190_sv2v_reg  <= w_data_i[93];
      \nz.mem_189_sv2v_reg  <= w_data_i[92];
      \nz.mem_188_sv2v_reg  <= w_data_i[91];
      \nz.mem_187_sv2v_reg  <= w_data_i[90];
      \nz.mem_186_sv2v_reg  <= w_data_i[89];
      \nz.mem_185_sv2v_reg  <= w_data_i[88];
      \nz.mem_184_sv2v_reg  <= w_data_i[87];
      \nz.mem_183_sv2v_reg  <= w_data_i[86];
      \nz.mem_182_sv2v_reg  <= w_data_i[85];
      \nz.mem_181_sv2v_reg  <= w_data_i[84];
      \nz.mem_180_sv2v_reg  <= w_data_i[83];
      \nz.mem_179_sv2v_reg  <= w_data_i[82];
      \nz.mem_178_sv2v_reg  <= w_data_i[81];
      \nz.mem_177_sv2v_reg  <= w_data_i[80];
      \nz.mem_176_sv2v_reg  <= w_data_i[79];
      \nz.mem_175_sv2v_reg  <= w_data_i[78];
      \nz.mem_174_sv2v_reg  <= w_data_i[77];
      \nz.mem_173_sv2v_reg  <= w_data_i[76];
      \nz.mem_172_sv2v_reg  <= w_data_i[75];
      \nz.mem_171_sv2v_reg  <= w_data_i[74];
      \nz.mem_170_sv2v_reg  <= w_data_i[73];
      \nz.mem_169_sv2v_reg  <= w_data_i[72];
      \nz.mem_168_sv2v_reg  <= w_data_i[71];
      \nz.mem_167_sv2v_reg  <= w_data_i[70];
      \nz.mem_166_sv2v_reg  <= w_data_i[69];
      \nz.mem_165_sv2v_reg  <= w_data_i[68];
      \nz.mem_164_sv2v_reg  <= w_data_i[67];
      \nz.mem_163_sv2v_reg  <= w_data_i[66];
      \nz.mem_162_sv2v_reg  <= w_data_i[65];
      \nz.mem_161_sv2v_reg  <= w_data_i[64];
      \nz.mem_160_sv2v_reg  <= w_data_i[63];
      \nz.mem_159_sv2v_reg  <= w_data_i[62];
      \nz.mem_158_sv2v_reg  <= w_data_i[61];
      \nz.mem_157_sv2v_reg  <= w_data_i[60];
      \nz.mem_156_sv2v_reg  <= w_data_i[59];
      \nz.mem_155_sv2v_reg  <= w_data_i[58];
      \nz.mem_154_sv2v_reg  <= w_data_i[57];
      \nz.mem_153_sv2v_reg  <= w_data_i[56];
      \nz.mem_152_sv2v_reg  <= w_data_i[55];
      \nz.mem_151_sv2v_reg  <= w_data_i[54];
      \nz.mem_150_sv2v_reg  <= w_data_i[53];
      \nz.mem_149_sv2v_reg  <= w_data_i[52];
      \nz.mem_148_sv2v_reg  <= w_data_i[51];
      \nz.mem_147_sv2v_reg  <= w_data_i[50];
      \nz.mem_146_sv2v_reg  <= w_data_i[49];
      \nz.mem_145_sv2v_reg  <= w_data_i[48];
      \nz.mem_144_sv2v_reg  <= w_data_i[47];
      \nz.mem_143_sv2v_reg  <= w_data_i[46];
      \nz.mem_142_sv2v_reg  <= w_data_i[45];
      \nz.mem_141_sv2v_reg  <= w_data_i[44];
      \nz.mem_140_sv2v_reg  <= w_data_i[43];
      \nz.mem_139_sv2v_reg  <= w_data_i[42];
      \nz.mem_138_sv2v_reg  <= w_data_i[41];
      \nz.mem_137_sv2v_reg  <= w_data_i[40];
      \nz.mem_136_sv2v_reg  <= w_data_i[39];
      \nz.mem_135_sv2v_reg  <= w_data_i[38];
      \nz.mem_134_sv2v_reg  <= w_data_i[37];
      \nz.mem_133_sv2v_reg  <= w_data_i[36];
      \nz.mem_132_sv2v_reg  <= w_data_i[35];
      \nz.mem_131_sv2v_reg  <= w_data_i[34];
      \nz.mem_130_sv2v_reg  <= w_data_i[33];
      \nz.mem_129_sv2v_reg  <= w_data_i[32];
      \nz.mem_128_sv2v_reg  <= w_data_i[31];
      \nz.mem_127_sv2v_reg  <= w_data_i[30];
      \nz.mem_126_sv2v_reg  <= w_data_i[29];
      \nz.mem_125_sv2v_reg  <= w_data_i[28];
      \nz.mem_124_sv2v_reg  <= w_data_i[27];
      \nz.mem_123_sv2v_reg  <= w_data_i[26];
      \nz.mem_122_sv2v_reg  <= w_data_i[25];
      \nz.mem_121_sv2v_reg  <= w_data_i[24];
      \nz.mem_120_sv2v_reg  <= w_data_i[23];
      \nz.mem_119_sv2v_reg  <= w_data_i[22];
      \nz.mem_118_sv2v_reg  <= w_data_i[21];
      \nz.mem_117_sv2v_reg  <= w_data_i[20];
      \nz.mem_116_sv2v_reg  <= w_data_i[19];
      \nz.mem_115_sv2v_reg  <= w_data_i[18];
      \nz.mem_114_sv2v_reg  <= w_data_i[17];
      \nz.mem_113_sv2v_reg  <= w_data_i[16];
      \nz.mem_112_sv2v_reg  <= w_data_i[15];
      \nz.mem_111_sv2v_reg  <= w_data_i[14];
      \nz.mem_110_sv2v_reg  <= w_data_i[13];
      \nz.mem_109_sv2v_reg  <= w_data_i[12];
      \nz.mem_108_sv2v_reg  <= w_data_i[11];
      \nz.mem_107_sv2v_reg  <= w_data_i[10];
      \nz.mem_106_sv2v_reg  <= w_data_i[9];
      \nz.mem_105_sv2v_reg  <= w_data_i[8];
      \nz.mem_104_sv2v_reg  <= w_data_i[7];
      \nz.mem_103_sv2v_reg  <= w_data_i[6];
      \nz.mem_102_sv2v_reg  <= w_data_i[5];
      \nz.mem_101_sv2v_reg  <= w_data_i[4];
      \nz.mem_100_sv2v_reg  <= w_data_i[3];
      \nz.mem_99_sv2v_reg  <= w_data_i[2];
      \nz.mem_98_sv2v_reg  <= w_data_i[1];
      \nz.mem_97_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_96_sv2v_reg  <= w_data_i[96];
      \nz.mem_95_sv2v_reg  <= w_data_i[95];
      \nz.mem_94_sv2v_reg  <= w_data_i[94];
      \nz.mem_93_sv2v_reg  <= w_data_i[93];
      \nz.mem_92_sv2v_reg  <= w_data_i[92];
      \nz.mem_91_sv2v_reg  <= w_data_i[91];
      \nz.mem_90_sv2v_reg  <= w_data_i[90];
      \nz.mem_89_sv2v_reg  <= w_data_i[89];
      \nz.mem_88_sv2v_reg  <= w_data_i[88];
      \nz.mem_87_sv2v_reg  <= w_data_i[87];
      \nz.mem_86_sv2v_reg  <= w_data_i[86];
      \nz.mem_85_sv2v_reg  <= w_data_i[85];
      \nz.mem_84_sv2v_reg  <= w_data_i[84];
      \nz.mem_83_sv2v_reg  <= w_data_i[83];
      \nz.mem_82_sv2v_reg  <= w_data_i[82];
      \nz.mem_81_sv2v_reg  <= w_data_i[81];
      \nz.mem_80_sv2v_reg  <= w_data_i[80];
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p97_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [96:0] w_data_i;
  input [0:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;

  bsg_mem_1r1w_synth_width_p97_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p97_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [96:0] data_i;
  output [96:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [96:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p97_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_fifo_1r1w_small_width_p97_els_p2
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [96:0] data_i;
  output [96:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [96:0] data_o;
  wire ready_o,v_o;

  bsg_two_fifo_width_p97_ready_THEN_valid_p0
  \unhardened.tf.twof 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_i(v_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s01_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,y_gt,y_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign req_o[2] = x_dirs_i > my_x_i;
  assign y_gt = y_dirs_i > my_y_i;
  assign req_o[1] = N0 & N1;
  assign N0 = ~req_o[2];
  assign N1 = ~x_eq;
  assign y_lt = N2 & N3;
  assign N2 = ~y_gt;
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[3] = x_eq & y_lt;
  assign req_o[4] = x_eq & y_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s02_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,y_gt,y_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign req_o[2] = x_dirs_i > my_x_i;
  assign y_gt = y_dirs_i > my_y_i;
  assign req_o[1] = N0 & N1;
  assign N0 = ~req_o[2];
  assign N1 = ~x_eq;
  assign y_lt = N2 & N3;
  assign N2 = ~y_gt;
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[3] = x_eq & y_lt;
  assign req_o[4] = x_eq & y_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s04_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,y_gt,y_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign req_o[2] = x_dirs_i > my_x_i;
  assign y_gt = y_dirs_i > my_y_i;
  assign req_o[1] = N0 & N1;
  assign N0 = ~req_o[2];
  assign N1 = ~x_eq;
  assign y_lt = N2 & N3;
  assign N2 = ~y_gt;
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[3] = x_eq & y_lt;
  assign req_o[4] = x_eq & y_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s08_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,y_gt,y_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign req_o[2] = x_dirs_i > my_x_i;
  assign y_gt = y_dirs_i > my_y_i;
  assign req_o[1] = N0 & N1;
  assign N0 = ~req_o[2];
  assign N1 = ~x_eq;
  assign y_lt = N2 & N3;
  assign N2 = ~y_gt;
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[3] = x_eq & y_lt;
  assign req_o[4] = x_eq & y_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s10_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,y_gt,y_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign req_o[2] = x_dirs_i > my_x_i;
  assign y_gt = y_dirs_i > my_y_i;
  assign req_o[1] = N0 & N1;
  assign N0 = ~req_o[2];
  assign N1 = ~x_eq;
  assign y_lt = N2 & N3;
  assign N2 = ~y_gt;
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[3] = x_eq & y_lt;
  assign req_o[4] = x_eq & y_gt;

endmodule



module bsg_transpose_width_p5_els_p5
(
  i,
  o
);

  input [24:0] i;
  output [24:0] o;
  wire [24:0] o;
  assign o[24] = i[24];
  assign o[23] = i[19];
  assign o[22] = i[14];
  assign o[21] = i[9];
  assign o[20] = i[4];
  assign o[19] = i[23];
  assign o[18] = i[18];
  assign o[17] = i[13];
  assign o[16] = i[8];
  assign o[15] = i[3];
  assign o[14] = i[22];
  assign o[13] = i[17];
  assign o[12] = i[12];
  assign o[11] = i[7];
  assign o[10] = i[2];
  assign o[9] = i[21];
  assign o[8] = i[16];
  assign o[7] = i[11];
  assign o[6] = i[6];
  assign o[5] = i[1];
  assign o[4] = i[20];
  assign o[3] = i[15];
  assign o[2] = i[10];
  assign o[1] = i[5];
  assign o[0] = i[0];

endmodule



module bsg_array_concentrate_static_1f_97
(
  i,
  o
);

  input [484:0] i;
  output [484:0] o;
  wire [484:0] o;
  assign o[484] = i[484];
  assign o[483] = i[483];
  assign o[482] = i[482];
  assign o[481] = i[481];
  assign o[480] = i[480];
  assign o[479] = i[479];
  assign o[478] = i[478];
  assign o[477] = i[477];
  assign o[476] = i[476];
  assign o[475] = i[475];
  assign o[474] = i[474];
  assign o[473] = i[473];
  assign o[472] = i[472];
  assign o[471] = i[471];
  assign o[470] = i[470];
  assign o[469] = i[469];
  assign o[468] = i[468];
  assign o[467] = i[467];
  assign o[466] = i[466];
  assign o[465] = i[465];
  assign o[464] = i[464];
  assign o[463] = i[463];
  assign o[462] = i[462];
  assign o[461] = i[461];
  assign o[460] = i[460];
  assign o[459] = i[459];
  assign o[458] = i[458];
  assign o[457] = i[457];
  assign o[456] = i[456];
  assign o[455] = i[455];
  assign o[454] = i[454];
  assign o[453] = i[453];
  assign o[452] = i[452];
  assign o[451] = i[451];
  assign o[450] = i[450];
  assign o[449] = i[449];
  assign o[448] = i[448];
  assign o[447] = i[447];
  assign o[446] = i[446];
  assign o[445] = i[445];
  assign o[444] = i[444];
  assign o[443] = i[443];
  assign o[442] = i[442];
  assign o[441] = i[441];
  assign o[440] = i[440];
  assign o[439] = i[439];
  assign o[438] = i[438];
  assign o[437] = i[437];
  assign o[436] = i[436];
  assign o[435] = i[435];
  assign o[434] = i[434];
  assign o[433] = i[433];
  assign o[432] = i[432];
  assign o[431] = i[431];
  assign o[430] = i[430];
  assign o[429] = i[429];
  assign o[428] = i[428];
  assign o[427] = i[427];
  assign o[426] = i[426];
  assign o[425] = i[425];
  assign o[424] = i[424];
  assign o[423] = i[423];
  assign o[422] = i[422];
  assign o[421] = i[421];
  assign o[420] = i[420];
  assign o[419] = i[419];
  assign o[418] = i[418];
  assign o[417] = i[417];
  assign o[416] = i[416];
  assign o[415] = i[415];
  assign o[414] = i[414];
  assign o[413] = i[413];
  assign o[412] = i[412];
  assign o[411] = i[411];
  assign o[410] = i[410];
  assign o[409] = i[409];
  assign o[408] = i[408];
  assign o[407] = i[407];
  assign o[406] = i[406];
  assign o[405] = i[405];
  assign o[404] = i[404];
  assign o[403] = i[403];
  assign o[402] = i[402];
  assign o[401] = i[401];
  assign o[400] = i[400];
  assign o[399] = i[399];
  assign o[398] = i[398];
  assign o[397] = i[397];
  assign o[396] = i[396];
  assign o[395] = i[395];
  assign o[394] = i[394];
  assign o[393] = i[393];
  assign o[392] = i[392];
  assign o[391] = i[391];
  assign o[390] = i[390];
  assign o[389] = i[389];
  assign o[388] = i[388];
  assign o[387] = i[387];
  assign o[386] = i[386];
  assign o[385] = i[385];
  assign o[384] = i[384];
  assign o[383] = i[383];
  assign o[382] = i[382];
  assign o[381] = i[381];
  assign o[380] = i[380];
  assign o[379] = i[379];
  assign o[378] = i[378];
  assign o[377] = i[377];
  assign o[376] = i[376];
  assign o[375] = i[375];
  assign o[374] = i[374];
  assign o[373] = i[373];
  assign o[372] = i[372];
  assign o[371] = i[371];
  assign o[370] = i[370];
  assign o[369] = i[369];
  assign o[368] = i[368];
  assign o[367] = i[367];
  assign o[366] = i[366];
  assign o[365] = i[365];
  assign o[364] = i[364];
  assign o[363] = i[363];
  assign o[362] = i[362];
  assign o[361] = i[361];
  assign o[360] = i[360];
  assign o[359] = i[359];
  assign o[358] = i[358];
  assign o[357] = i[357];
  assign o[356] = i[356];
  assign o[355] = i[355];
  assign o[354] = i[354];
  assign o[353] = i[353];
  assign o[352] = i[352];
  assign o[351] = i[351];
  assign o[350] = i[350];
  assign o[349] = i[349];
  assign o[348] = i[348];
  assign o[347] = i[347];
  assign o[346] = i[346];
  assign o[345] = i[345];
  assign o[344] = i[344];
  assign o[343] = i[343];
  assign o[342] = i[342];
  assign o[341] = i[341];
  assign o[340] = i[340];
  assign o[339] = i[339];
  assign o[338] = i[338];
  assign o[337] = i[337];
  assign o[336] = i[336];
  assign o[335] = i[335];
  assign o[334] = i[334];
  assign o[333] = i[333];
  assign o[332] = i[332];
  assign o[331] = i[331];
  assign o[330] = i[330];
  assign o[329] = i[329];
  assign o[328] = i[328];
  assign o[327] = i[327];
  assign o[326] = i[326];
  assign o[325] = i[325];
  assign o[324] = i[324];
  assign o[323] = i[323];
  assign o[322] = i[322];
  assign o[321] = i[321];
  assign o[320] = i[320];
  assign o[319] = i[319];
  assign o[318] = i[318];
  assign o[317] = i[317];
  assign o[316] = i[316];
  assign o[315] = i[315];
  assign o[314] = i[314];
  assign o[313] = i[313];
  assign o[312] = i[312];
  assign o[311] = i[311];
  assign o[310] = i[310];
  assign o[309] = i[309];
  assign o[308] = i[308];
  assign o[307] = i[307];
  assign o[306] = i[306];
  assign o[305] = i[305];
  assign o[304] = i[304];
  assign o[303] = i[303];
  assign o[302] = i[302];
  assign o[301] = i[301];
  assign o[300] = i[300];
  assign o[299] = i[299];
  assign o[298] = i[298];
  assign o[297] = i[297];
  assign o[296] = i[296];
  assign o[295] = i[295];
  assign o[294] = i[294];
  assign o[293] = i[293];
  assign o[292] = i[292];
  assign o[291] = i[291];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_1f
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_scan_0000000a_1
(
  i,
  o
);

  input [9:0] i;
  output [9:0] o;
  wire [9:0] o;
  wire t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,
  t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,
  t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__9_ = i[9] | 1'b0;
  assign t_1__8_ = i[8] | i[9];
  assign t_1__7_ = i[7] | i[8];
  assign t_1__6_ = i[6] | i[7];
  assign t_1__5_ = i[5] | i[6];
  assign t_1__4_ = i[4] | i[5];
  assign t_1__3_ = i[3] | i[4];
  assign t_1__2_ = i[2] | i[3];
  assign t_1__1_ = i[1] | i[2];
  assign t_1__0_ = i[0] | i[1];
  assign t_2__9_ = t_1__9_ | 1'b0;
  assign t_2__8_ = t_1__8_ | 1'b0;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__9_ = t_2__9_ | 1'b0;
  assign t_3__8_ = t_2__8_ | 1'b0;
  assign t_3__7_ = t_2__7_ | 1'b0;
  assign t_3__6_ = t_2__6_ | 1'b0;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign o[9] = t_3__9_ | 1'b0;
  assign o[8] = t_3__8_ | 1'b0;
  assign o[7] = t_3__7_ | 1'b0;
  assign o[6] = t_3__6_ | 1'b0;
  assign o[5] = t_3__5_ | 1'b0;
  assign o[4] = t_3__4_ | 1'b0;
  assign o[3] = t_3__3_ | 1'b0;
  assign o[2] = t_3__2_ | 1'b0;
  assign o[1] = t_3__1_ | t_3__9_;
  assign o[0] = t_3__0_ | t_3__8_;

endmodule



module bsg_arb_round_robin_05
(
  clk_i,
  reset_i,
  reqs_i,
  grants_o,
  yumi_i
);

  input [4:0] reqs_i;
  output [4:0] grants_o;
  input clk_i;
  input reset_i;
  input yumi_i;
  wire [4:0] grants_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;
  wire [3:0] \fi2.thermocode_r ,\fi2.thermocode_n ;
  wire [8:5] \fi2.scan_li ;
  wire [9:0] \fi2.scan_lo ;
  wire [8:0] \fi2.edge_detect ;
  reg \fi2.thermocode_r_3_sv2v_reg ,\fi2.thermocode_r_2_sv2v_reg ,
  \fi2.thermocode_r_1_sv2v_reg ,\fi2.thermocode_r_0_sv2v_reg ;
  assign \fi2.thermocode_r [3] = \fi2.thermocode_r_3_sv2v_reg ;
  assign \fi2.thermocode_r [2] = \fi2.thermocode_r_2_sv2v_reg ;
  assign \fi2.thermocode_r [1] = \fi2.thermocode_r_1_sv2v_reg ;
  assign \fi2.thermocode_r [0] = \fi2.thermocode_r_0_sv2v_reg ;

  bsg_scan_0000000a_1
  \fi2.scan 
  (
    .i({ 1'b0, \fi2.scan_li , reqs_i }),
    .o(\fi2.scan_lo )
  );

  assign N3 = (N0)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = yumi_i;
  assign \fi2.thermocode_n  = (N1)? \fi2.scan_lo [9:6] : 
                              (N5)? \fi2.scan_lo [4:1] : 1'b0;
  assign N1 = N4;
  assign N2 = ~yumi_i;
  assign \fi2.scan_li [8] = \fi2.thermocode_r [3] & reqs_i[3];
  assign \fi2.scan_li [7] = \fi2.thermocode_r [2] & reqs_i[2];
  assign \fi2.scan_li [6] = \fi2.thermocode_r [1] & reqs_i[1];
  assign \fi2.scan_li [5] = \fi2.thermocode_r [0] & reqs_i[0];
  assign \fi2.edge_detect [8] = N6 & \fi2.scan_lo [8];
  assign N6 = ~\fi2.scan_lo [9];
  assign \fi2.edge_detect [7] = N7 & \fi2.scan_lo [7];
  assign N7 = ~\fi2.scan_lo [8];
  assign \fi2.edge_detect [6] = N8 & \fi2.scan_lo [6];
  assign N8 = ~\fi2.scan_lo [7];
  assign \fi2.edge_detect [5] = N9 & \fi2.scan_lo [5];
  assign N9 = ~\fi2.scan_lo [6];
  assign \fi2.edge_detect [4] = N10 & \fi2.scan_lo [4];
  assign N10 = ~\fi2.scan_lo [5];
  assign \fi2.edge_detect [3] = N11 & \fi2.scan_lo [3];
  assign N11 = ~\fi2.scan_lo [4];
  assign \fi2.edge_detect [2] = N12 & \fi2.scan_lo [2];
  assign N12 = ~\fi2.scan_lo [3];
  assign \fi2.edge_detect [1] = N13 & \fi2.scan_lo [1];
  assign N13 = ~\fi2.scan_lo [2];
  assign \fi2.edge_detect [0] = N14 & \fi2.scan_lo [0];
  assign N14 = ~\fi2.scan_lo [1];
  assign grants_o[4] = \fi2.scan_lo [9] | \fi2.edge_detect [4];
  assign grants_o[3] = \fi2.edge_detect [8] | \fi2.edge_detect [3];
  assign grants_o[2] = \fi2.edge_detect [7] | \fi2.edge_detect [2];
  assign grants_o[1] = \fi2.edge_detect [6] | \fi2.edge_detect [1];
  assign grants_o[0] = \fi2.edge_detect [5] | \fi2.edge_detect [0];
  assign N4 = N17 | \fi2.scan_li [5];
  assign N17 = N16 | \fi2.scan_li [6];
  assign N16 = N15 | \fi2.scan_li [7];
  assign N15 = 1'b0 | \fi2.scan_li [8];
  assign N5 = ~N4;

  always @(posedge clk_i) begin
    if(reset_i) begin
      \fi2.thermocode_r_3_sv2v_reg  <= 1'b0;
      \fi2.thermocode_r_2_sv2v_reg  <= 1'b0;
      \fi2.thermocode_r_1_sv2v_reg  <= 1'b0;
      \fi2.thermocode_r_0_sv2v_reg  <= 1'b0;
    end else if(N3) begin
      \fi2.thermocode_r_3_sv2v_reg  <= \fi2.thermocode_n [3];
      \fi2.thermocode_r_2_sv2v_reg  <= \fi2.thermocode_n [2];
      \fi2.thermocode_r_1_sv2v_reg  <= \fi2.thermocode_n [1];
      \fi2.thermocode_r_0_sv2v_reg  <= \fi2.thermocode_n [0];
    end 
  end


endmodule



module bsg_mux_one_hot_97_05
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [484:0] data_i;
  input [4:0] sel_one_hot_i;
  output [96:0] data_o;
  wire [96:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290;
  wire [484:0] data_masked;
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[2];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[2];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[2];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[2];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[2];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[2];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[2];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[2];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[2];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[2];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[2];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[2];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[2];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[2];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[2];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[2];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[2];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[2];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[2];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[2];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[2];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[2];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[2];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[2];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[2];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[2];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[2];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[2];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[2];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[2];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[2];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[2];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[2];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[2];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[2];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[2];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[2];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[2];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[2];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[2];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[2];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[2];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[2];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[2];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[2];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[2];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[2];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[2];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[2];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[2];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[2];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[2];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[2];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[2];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[2];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[2];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[2];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[2];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[2];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[2];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[2];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[2];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[2];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[2];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[2];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[2];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[3];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[3];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[3];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[3];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[3];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[3];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[3];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[3];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[3];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[3];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[3];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[3];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[3];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[3];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[3];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[3];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[3];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[3];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[3];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[3];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[3];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[3];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[3];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[3];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[3];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[3];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[3];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[3];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[3];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[3];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[3];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[3];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[3];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[3];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[3];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[3];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[3];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[3];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[3];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[3];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[3];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[3];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[3];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[3];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[3];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[3];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[3];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[3];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[3];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[3];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[3];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[3];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[3];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[3];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[3];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[3];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[3];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[3];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[3];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[3];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[3];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[3];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[3];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[3];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[3];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[3];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[3];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[3];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[3];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[3];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[3];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[3];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[3];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[3];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[3];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[3];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[3];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[3];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[3];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[3];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[3];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[3];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[3];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[3];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[3];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[3];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[3];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[3];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[3];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[3];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[3];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[3];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[3];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[3];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[3];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[4];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[4];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[4];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[4];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[4];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[4];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[4];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[4];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[4];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[4];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[4];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[4];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[4];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[4];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[4];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[4];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[4];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[4];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[4];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[4];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[4];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[4];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[4];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[4];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[4];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[4];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[4];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[4];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[4];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[4];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[4];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[4];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[4];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[4];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[4];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[4];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[4];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[4];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[4];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[4];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[4];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[4];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[4];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[4];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[4];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[4];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[4];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[4];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[4];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[4];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[4];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[4];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[4];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[4];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[4];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[4];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[4];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[4];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[4];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[4];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[4];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[4];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[4];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[4];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[4];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[4];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[4];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[4];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[4];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[4];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[4];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[4];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[4];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[4];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[4];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[4];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[4];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[4];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[4];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[4];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[4];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[4];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[4];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[4];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[4];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[4];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[4];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[4];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[4];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[4];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[4];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[4];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[4];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[4];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[4];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[4];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[97];
  assign N1 = N0 | data_masked[194];
  assign N0 = data_masked[388] | data_masked[291];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[98];
  assign N4 = N3 | data_masked[195];
  assign N3 = data_masked[389] | data_masked[292];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[99];
  assign N7 = N6 | data_masked[196];
  assign N6 = data_masked[390] | data_masked[293];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[100];
  assign N10 = N9 | data_masked[197];
  assign N9 = data_masked[391] | data_masked[294];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[101];
  assign N13 = N12 | data_masked[198];
  assign N12 = data_masked[392] | data_masked[295];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[102];
  assign N16 = N15 | data_masked[199];
  assign N15 = data_masked[393] | data_masked[296];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[103];
  assign N19 = N18 | data_masked[200];
  assign N18 = data_masked[394] | data_masked[297];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[104];
  assign N22 = N21 | data_masked[201];
  assign N21 = data_masked[395] | data_masked[298];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[105];
  assign N25 = N24 | data_masked[202];
  assign N24 = data_masked[396] | data_masked[299];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[106];
  assign N28 = N27 | data_masked[203];
  assign N27 = data_masked[397] | data_masked[300];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[107];
  assign N31 = N30 | data_masked[204];
  assign N30 = data_masked[398] | data_masked[301];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[108];
  assign N34 = N33 | data_masked[205];
  assign N33 = data_masked[399] | data_masked[302];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[109];
  assign N37 = N36 | data_masked[206];
  assign N36 = data_masked[400] | data_masked[303];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[110];
  assign N40 = N39 | data_masked[207];
  assign N39 = data_masked[401] | data_masked[304];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[111];
  assign N43 = N42 | data_masked[208];
  assign N42 = data_masked[402] | data_masked[305];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[112];
  assign N46 = N45 | data_masked[209];
  assign N45 = data_masked[403] | data_masked[306];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[113];
  assign N49 = N48 | data_masked[210];
  assign N48 = data_masked[404] | data_masked[307];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[114];
  assign N52 = N51 | data_masked[211];
  assign N51 = data_masked[405] | data_masked[308];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[115];
  assign N55 = N54 | data_masked[212];
  assign N54 = data_masked[406] | data_masked[309];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[116];
  assign N58 = N57 | data_masked[213];
  assign N57 = data_masked[407] | data_masked[310];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[117];
  assign N61 = N60 | data_masked[214];
  assign N60 = data_masked[408] | data_masked[311];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[118];
  assign N64 = N63 | data_masked[215];
  assign N63 = data_masked[409] | data_masked[312];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[119];
  assign N67 = N66 | data_masked[216];
  assign N66 = data_masked[410] | data_masked[313];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[120];
  assign N70 = N69 | data_masked[217];
  assign N69 = data_masked[411] | data_masked[314];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[121];
  assign N73 = N72 | data_masked[218];
  assign N72 = data_masked[412] | data_masked[315];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[122];
  assign N76 = N75 | data_masked[219];
  assign N75 = data_masked[413] | data_masked[316];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[123];
  assign N79 = N78 | data_masked[220];
  assign N78 = data_masked[414] | data_masked[317];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[124];
  assign N82 = N81 | data_masked[221];
  assign N81 = data_masked[415] | data_masked[318];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[125];
  assign N85 = N84 | data_masked[222];
  assign N84 = data_masked[416] | data_masked[319];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[126];
  assign N88 = N87 | data_masked[223];
  assign N87 = data_masked[417] | data_masked[320];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[127];
  assign N91 = N90 | data_masked[224];
  assign N90 = data_masked[418] | data_masked[321];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[128];
  assign N94 = N93 | data_masked[225];
  assign N93 = data_masked[419] | data_masked[322];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[129];
  assign N97 = N96 | data_masked[226];
  assign N96 = data_masked[420] | data_masked[323];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[130];
  assign N100 = N99 | data_masked[227];
  assign N99 = data_masked[421] | data_masked[324];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[131];
  assign N103 = N102 | data_masked[228];
  assign N102 = data_masked[422] | data_masked[325];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[132];
  assign N106 = N105 | data_masked[229];
  assign N105 = data_masked[423] | data_masked[326];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[133];
  assign N109 = N108 | data_masked[230];
  assign N108 = data_masked[424] | data_masked[327];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[134];
  assign N112 = N111 | data_masked[231];
  assign N111 = data_masked[425] | data_masked[328];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[135];
  assign N115 = N114 | data_masked[232];
  assign N114 = data_masked[426] | data_masked[329];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[136];
  assign N118 = N117 | data_masked[233];
  assign N117 = data_masked[427] | data_masked[330];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[137];
  assign N121 = N120 | data_masked[234];
  assign N120 = data_masked[428] | data_masked[331];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[138];
  assign N124 = N123 | data_masked[235];
  assign N123 = data_masked[429] | data_masked[332];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[139];
  assign N127 = N126 | data_masked[236];
  assign N126 = data_masked[430] | data_masked[333];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[140];
  assign N130 = N129 | data_masked[237];
  assign N129 = data_masked[431] | data_masked[334];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[141];
  assign N133 = N132 | data_masked[238];
  assign N132 = data_masked[432] | data_masked[335];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[142];
  assign N136 = N135 | data_masked[239];
  assign N135 = data_masked[433] | data_masked[336];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[143];
  assign N139 = N138 | data_masked[240];
  assign N138 = data_masked[434] | data_masked[337];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[144];
  assign N142 = N141 | data_masked[241];
  assign N141 = data_masked[435] | data_masked[338];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[145];
  assign N145 = N144 | data_masked[242];
  assign N144 = data_masked[436] | data_masked[339];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[146];
  assign N148 = N147 | data_masked[243];
  assign N147 = data_masked[437] | data_masked[340];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[147];
  assign N151 = N150 | data_masked[244];
  assign N150 = data_masked[438] | data_masked[341];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[148];
  assign N154 = N153 | data_masked[245];
  assign N153 = data_masked[439] | data_masked[342];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[149];
  assign N157 = N156 | data_masked[246];
  assign N156 = data_masked[440] | data_masked[343];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[150];
  assign N160 = N159 | data_masked[247];
  assign N159 = data_masked[441] | data_masked[344];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[151];
  assign N163 = N162 | data_masked[248];
  assign N162 = data_masked[442] | data_masked[345];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[152];
  assign N166 = N165 | data_masked[249];
  assign N165 = data_masked[443] | data_masked[346];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[153];
  assign N169 = N168 | data_masked[250];
  assign N168 = data_masked[444] | data_masked[347];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[154];
  assign N172 = N171 | data_masked[251];
  assign N171 = data_masked[445] | data_masked[348];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[155];
  assign N175 = N174 | data_masked[252];
  assign N174 = data_masked[446] | data_masked[349];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[156];
  assign N178 = N177 | data_masked[253];
  assign N177 = data_masked[447] | data_masked[350];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[157];
  assign N181 = N180 | data_masked[254];
  assign N180 = data_masked[448] | data_masked[351];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[158];
  assign N184 = N183 | data_masked[255];
  assign N183 = data_masked[449] | data_masked[352];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[159];
  assign N187 = N186 | data_masked[256];
  assign N186 = data_masked[450] | data_masked[353];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[160];
  assign N190 = N189 | data_masked[257];
  assign N189 = data_masked[451] | data_masked[354];
  assign data_o[64] = N194 | data_masked[64];
  assign N194 = N193 | data_masked[161];
  assign N193 = N192 | data_masked[258];
  assign N192 = data_masked[452] | data_masked[355];
  assign data_o[65] = N197 | data_masked[65];
  assign N197 = N196 | data_masked[162];
  assign N196 = N195 | data_masked[259];
  assign N195 = data_masked[453] | data_masked[356];
  assign data_o[66] = N200 | data_masked[66];
  assign N200 = N199 | data_masked[163];
  assign N199 = N198 | data_masked[260];
  assign N198 = data_masked[454] | data_masked[357];
  assign data_o[67] = N203 | data_masked[67];
  assign N203 = N202 | data_masked[164];
  assign N202 = N201 | data_masked[261];
  assign N201 = data_masked[455] | data_masked[358];
  assign data_o[68] = N206 | data_masked[68];
  assign N206 = N205 | data_masked[165];
  assign N205 = N204 | data_masked[262];
  assign N204 = data_masked[456] | data_masked[359];
  assign data_o[69] = N209 | data_masked[69];
  assign N209 = N208 | data_masked[166];
  assign N208 = N207 | data_masked[263];
  assign N207 = data_masked[457] | data_masked[360];
  assign data_o[70] = N212 | data_masked[70];
  assign N212 = N211 | data_masked[167];
  assign N211 = N210 | data_masked[264];
  assign N210 = data_masked[458] | data_masked[361];
  assign data_o[71] = N215 | data_masked[71];
  assign N215 = N214 | data_masked[168];
  assign N214 = N213 | data_masked[265];
  assign N213 = data_masked[459] | data_masked[362];
  assign data_o[72] = N218 | data_masked[72];
  assign N218 = N217 | data_masked[169];
  assign N217 = N216 | data_masked[266];
  assign N216 = data_masked[460] | data_masked[363];
  assign data_o[73] = N221 | data_masked[73];
  assign N221 = N220 | data_masked[170];
  assign N220 = N219 | data_masked[267];
  assign N219 = data_masked[461] | data_masked[364];
  assign data_o[74] = N224 | data_masked[74];
  assign N224 = N223 | data_masked[171];
  assign N223 = N222 | data_masked[268];
  assign N222 = data_masked[462] | data_masked[365];
  assign data_o[75] = N227 | data_masked[75];
  assign N227 = N226 | data_masked[172];
  assign N226 = N225 | data_masked[269];
  assign N225 = data_masked[463] | data_masked[366];
  assign data_o[76] = N230 | data_masked[76];
  assign N230 = N229 | data_masked[173];
  assign N229 = N228 | data_masked[270];
  assign N228 = data_masked[464] | data_masked[367];
  assign data_o[77] = N233 | data_masked[77];
  assign N233 = N232 | data_masked[174];
  assign N232 = N231 | data_masked[271];
  assign N231 = data_masked[465] | data_masked[368];
  assign data_o[78] = N236 | data_masked[78];
  assign N236 = N235 | data_masked[175];
  assign N235 = N234 | data_masked[272];
  assign N234 = data_masked[466] | data_masked[369];
  assign data_o[79] = N239 | data_masked[79];
  assign N239 = N238 | data_masked[176];
  assign N238 = N237 | data_masked[273];
  assign N237 = data_masked[467] | data_masked[370];
  assign data_o[80] = N242 | data_masked[80];
  assign N242 = N241 | data_masked[177];
  assign N241 = N240 | data_masked[274];
  assign N240 = data_masked[468] | data_masked[371];
  assign data_o[81] = N245 | data_masked[81];
  assign N245 = N244 | data_masked[178];
  assign N244 = N243 | data_masked[275];
  assign N243 = data_masked[469] | data_masked[372];
  assign data_o[82] = N248 | data_masked[82];
  assign N248 = N247 | data_masked[179];
  assign N247 = N246 | data_masked[276];
  assign N246 = data_masked[470] | data_masked[373];
  assign data_o[83] = N251 | data_masked[83];
  assign N251 = N250 | data_masked[180];
  assign N250 = N249 | data_masked[277];
  assign N249 = data_masked[471] | data_masked[374];
  assign data_o[84] = N254 | data_masked[84];
  assign N254 = N253 | data_masked[181];
  assign N253 = N252 | data_masked[278];
  assign N252 = data_masked[472] | data_masked[375];
  assign data_o[85] = N257 | data_masked[85];
  assign N257 = N256 | data_masked[182];
  assign N256 = N255 | data_masked[279];
  assign N255 = data_masked[473] | data_masked[376];
  assign data_o[86] = N260 | data_masked[86];
  assign N260 = N259 | data_masked[183];
  assign N259 = N258 | data_masked[280];
  assign N258 = data_masked[474] | data_masked[377];
  assign data_o[87] = N263 | data_masked[87];
  assign N263 = N262 | data_masked[184];
  assign N262 = N261 | data_masked[281];
  assign N261 = data_masked[475] | data_masked[378];
  assign data_o[88] = N266 | data_masked[88];
  assign N266 = N265 | data_masked[185];
  assign N265 = N264 | data_masked[282];
  assign N264 = data_masked[476] | data_masked[379];
  assign data_o[89] = N269 | data_masked[89];
  assign N269 = N268 | data_masked[186];
  assign N268 = N267 | data_masked[283];
  assign N267 = data_masked[477] | data_masked[380];
  assign data_o[90] = N272 | data_masked[90];
  assign N272 = N271 | data_masked[187];
  assign N271 = N270 | data_masked[284];
  assign N270 = data_masked[478] | data_masked[381];
  assign data_o[91] = N275 | data_masked[91];
  assign N275 = N274 | data_masked[188];
  assign N274 = N273 | data_masked[285];
  assign N273 = data_masked[479] | data_masked[382];
  assign data_o[92] = N278 | data_masked[92];
  assign N278 = N277 | data_masked[189];
  assign N277 = N276 | data_masked[286];
  assign N276 = data_masked[480] | data_masked[383];
  assign data_o[93] = N281 | data_masked[93];
  assign N281 = N280 | data_masked[190];
  assign N280 = N279 | data_masked[287];
  assign N279 = data_masked[481] | data_masked[384];
  assign data_o[94] = N284 | data_masked[94];
  assign N284 = N283 | data_masked[191];
  assign N283 = N282 | data_masked[288];
  assign N282 = data_masked[482] | data_masked[385];
  assign data_o[95] = N287 | data_masked[95];
  assign N287 = N286 | data_masked[192];
  assign N286 = N285 | data_masked[289];
  assign N285 = data_masked[483] | data_masked[386];
  assign data_o[96] = N290 | data_masked[96];
  assign N290 = N289 | data_masked[193];
  assign N289 = N288 | data_masked[290];
  assign N288 = data_masked[484] | data_masked[387];

endmodule



module bsg_unconcentrate_static_1f_0
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_array_concentrate_static_05_97
(
  i,
  o
);

  input [484:0] i;
  output [193:0] o;
  wire [193:0] o;
  assign o[193] = i[290];
  assign o[192] = i[289];
  assign o[191] = i[288];
  assign o[190] = i[287];
  assign o[189] = i[286];
  assign o[188] = i[285];
  assign o[187] = i[284];
  assign o[186] = i[283];
  assign o[185] = i[282];
  assign o[184] = i[281];
  assign o[183] = i[280];
  assign o[182] = i[279];
  assign o[181] = i[278];
  assign o[180] = i[277];
  assign o[179] = i[276];
  assign o[178] = i[275];
  assign o[177] = i[274];
  assign o[176] = i[273];
  assign o[175] = i[272];
  assign o[174] = i[271];
  assign o[173] = i[270];
  assign o[172] = i[269];
  assign o[171] = i[268];
  assign o[170] = i[267];
  assign o[169] = i[266];
  assign o[168] = i[265];
  assign o[167] = i[264];
  assign o[166] = i[263];
  assign o[165] = i[262];
  assign o[164] = i[261];
  assign o[163] = i[260];
  assign o[162] = i[259];
  assign o[161] = i[258];
  assign o[160] = i[257];
  assign o[159] = i[256];
  assign o[158] = i[255];
  assign o[157] = i[254];
  assign o[156] = i[253];
  assign o[155] = i[252];
  assign o[154] = i[251];
  assign o[153] = i[250];
  assign o[152] = i[249];
  assign o[151] = i[248];
  assign o[150] = i[247];
  assign o[149] = i[246];
  assign o[148] = i[245];
  assign o[147] = i[244];
  assign o[146] = i[243];
  assign o[145] = i[242];
  assign o[144] = i[241];
  assign o[143] = i[240];
  assign o[142] = i[239];
  assign o[141] = i[238];
  assign o[140] = i[237];
  assign o[139] = i[236];
  assign o[138] = i[235];
  assign o[137] = i[234];
  assign o[136] = i[233];
  assign o[135] = i[232];
  assign o[134] = i[231];
  assign o[133] = i[230];
  assign o[132] = i[229];
  assign o[131] = i[228];
  assign o[130] = i[227];
  assign o[129] = i[226];
  assign o[128] = i[225];
  assign o[127] = i[224];
  assign o[126] = i[223];
  assign o[125] = i[222];
  assign o[124] = i[221];
  assign o[123] = i[220];
  assign o[122] = i[219];
  assign o[121] = i[218];
  assign o[120] = i[217];
  assign o[119] = i[216];
  assign o[118] = i[215];
  assign o[117] = i[214];
  assign o[116] = i[213];
  assign o[115] = i[212];
  assign o[114] = i[211];
  assign o[113] = i[210];
  assign o[112] = i[209];
  assign o[111] = i[208];
  assign o[110] = i[207];
  assign o[109] = i[206];
  assign o[108] = i[205];
  assign o[107] = i[204];
  assign o[106] = i[203];
  assign o[105] = i[202];
  assign o[104] = i[201];
  assign o[103] = i[200];
  assign o[102] = i[199];
  assign o[101] = i[198];
  assign o[100] = i[197];
  assign o[99] = i[196];
  assign o[98] = i[195];
  assign o[97] = i[194];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_05
(
  i,
  o
);

  input [4:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[1] = i[2];
  assign o[0] = i[0];

endmodule



module bsg_scan_00000004_1
(
  i,
  o
);

  input [3:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__3_ = i[3] | 1'b0;
  assign t_1__2_ = i[2] | i[3];
  assign t_1__1_ = i[1] | i[2];
  assign t_1__0_ = i[0] | i[1];
  assign o[3] = t_1__3_ | 1'b0;
  assign o[2] = t_1__2_ | 1'b0;
  assign o[1] = t_1__1_ | t_1__3_;
  assign o[0] = t_1__0_ | t_1__2_;

endmodule



module bsg_arb_round_robin_02
(
  clk_i,
  reset_i,
  reqs_i,
  grants_o,
  yumi_i
);

  input [1:0] reqs_i;
  output [1:0] grants_o;
  input clk_i;
  input reset_i;
  input yumi_i;
  wire [1:0] grants_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8;
  wire [0:0] \fi2.thermocode_r ,\fi2.thermocode_n ;
  wire [2:2] \fi2.scan_li ;
  wire [3:0] \fi2.scan_lo ;
  wire [2:0] \fi2.edge_detect ;
  reg \fi2.thermocode_r_0_sv2v_reg ;
  assign \fi2.thermocode_r [0] = \fi2.thermocode_r_0_sv2v_reg ;

  bsg_scan_00000004_1
  \fi2.scan 
  (
    .i({ 1'b0, \fi2.scan_li [2:2], reqs_i }),
    .o(\fi2.scan_lo )
  );

  assign N3 = (N0)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = yumi_i;
  assign \fi2.thermocode_n [0] = (N1)? \fi2.scan_lo [3] : 
                                 (N5)? \fi2.scan_lo [1] : 1'b0;
  assign N1 = N4;
  assign N2 = ~yumi_i;
  assign \fi2.scan_li [2] = \fi2.thermocode_r [0] & reqs_i[0];
  assign \fi2.edge_detect [2] = N6 & \fi2.scan_lo [2];
  assign N6 = ~\fi2.scan_lo [3];
  assign \fi2.edge_detect [1] = N7 & \fi2.scan_lo [1];
  assign N7 = ~\fi2.scan_lo [2];
  assign \fi2.edge_detect [0] = N8 & \fi2.scan_lo [0];
  assign N8 = ~\fi2.scan_lo [1];
  assign grants_o[1] = \fi2.scan_lo [3] | \fi2.edge_detect [1];
  assign grants_o[0] = \fi2.edge_detect [2] | \fi2.edge_detect [0];
  assign N4 = 1'b0 | \fi2.scan_li [2];
  assign N5 = ~N4;

  always @(posedge clk_i) begin
    if(reset_i) begin
      \fi2.thermocode_r_0_sv2v_reg  <= 1'b0;
    end else if(N3) begin
      \fi2.thermocode_r_0_sv2v_reg  <= \fi2.thermocode_n [0];
    end 
  end


endmodule



module bsg_mux_one_hot_97_02
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [193:0] data_i;
  input [1:0] sel_one_hot_i;
  output [96:0] data_o;
  wire [96:0] data_o;
  wire [193:0] data_masked;
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[97] | data_masked[0];
  assign data_o[1] = data_masked[98] | data_masked[1];
  assign data_o[2] = data_masked[99] | data_masked[2];
  assign data_o[3] = data_masked[100] | data_masked[3];
  assign data_o[4] = data_masked[101] | data_masked[4];
  assign data_o[5] = data_masked[102] | data_masked[5];
  assign data_o[6] = data_masked[103] | data_masked[6];
  assign data_o[7] = data_masked[104] | data_masked[7];
  assign data_o[8] = data_masked[105] | data_masked[8];
  assign data_o[9] = data_masked[106] | data_masked[9];
  assign data_o[10] = data_masked[107] | data_masked[10];
  assign data_o[11] = data_masked[108] | data_masked[11];
  assign data_o[12] = data_masked[109] | data_masked[12];
  assign data_o[13] = data_masked[110] | data_masked[13];
  assign data_o[14] = data_masked[111] | data_masked[14];
  assign data_o[15] = data_masked[112] | data_masked[15];
  assign data_o[16] = data_masked[113] | data_masked[16];
  assign data_o[17] = data_masked[114] | data_masked[17];
  assign data_o[18] = data_masked[115] | data_masked[18];
  assign data_o[19] = data_masked[116] | data_masked[19];
  assign data_o[20] = data_masked[117] | data_masked[20];
  assign data_o[21] = data_masked[118] | data_masked[21];
  assign data_o[22] = data_masked[119] | data_masked[22];
  assign data_o[23] = data_masked[120] | data_masked[23];
  assign data_o[24] = data_masked[121] | data_masked[24];
  assign data_o[25] = data_masked[122] | data_masked[25];
  assign data_o[26] = data_masked[123] | data_masked[26];
  assign data_o[27] = data_masked[124] | data_masked[27];
  assign data_o[28] = data_masked[125] | data_masked[28];
  assign data_o[29] = data_masked[126] | data_masked[29];
  assign data_o[30] = data_masked[127] | data_masked[30];
  assign data_o[31] = data_masked[128] | data_masked[31];
  assign data_o[32] = data_masked[129] | data_masked[32];
  assign data_o[33] = data_masked[130] | data_masked[33];
  assign data_o[34] = data_masked[131] | data_masked[34];
  assign data_o[35] = data_masked[132] | data_masked[35];
  assign data_o[36] = data_masked[133] | data_masked[36];
  assign data_o[37] = data_masked[134] | data_masked[37];
  assign data_o[38] = data_masked[135] | data_masked[38];
  assign data_o[39] = data_masked[136] | data_masked[39];
  assign data_o[40] = data_masked[137] | data_masked[40];
  assign data_o[41] = data_masked[138] | data_masked[41];
  assign data_o[42] = data_masked[139] | data_masked[42];
  assign data_o[43] = data_masked[140] | data_masked[43];
  assign data_o[44] = data_masked[141] | data_masked[44];
  assign data_o[45] = data_masked[142] | data_masked[45];
  assign data_o[46] = data_masked[143] | data_masked[46];
  assign data_o[47] = data_masked[144] | data_masked[47];
  assign data_o[48] = data_masked[145] | data_masked[48];
  assign data_o[49] = data_masked[146] | data_masked[49];
  assign data_o[50] = data_masked[147] | data_masked[50];
  assign data_o[51] = data_masked[148] | data_masked[51];
  assign data_o[52] = data_masked[149] | data_masked[52];
  assign data_o[53] = data_masked[150] | data_masked[53];
  assign data_o[54] = data_masked[151] | data_masked[54];
  assign data_o[55] = data_masked[152] | data_masked[55];
  assign data_o[56] = data_masked[153] | data_masked[56];
  assign data_o[57] = data_masked[154] | data_masked[57];
  assign data_o[58] = data_masked[155] | data_masked[58];
  assign data_o[59] = data_masked[156] | data_masked[59];
  assign data_o[60] = data_masked[157] | data_masked[60];
  assign data_o[61] = data_masked[158] | data_masked[61];
  assign data_o[62] = data_masked[159] | data_masked[62];
  assign data_o[63] = data_masked[160] | data_masked[63];
  assign data_o[64] = data_masked[161] | data_masked[64];
  assign data_o[65] = data_masked[162] | data_masked[65];
  assign data_o[66] = data_masked[163] | data_masked[66];
  assign data_o[67] = data_masked[164] | data_masked[67];
  assign data_o[68] = data_masked[165] | data_masked[68];
  assign data_o[69] = data_masked[166] | data_masked[69];
  assign data_o[70] = data_masked[167] | data_masked[70];
  assign data_o[71] = data_masked[168] | data_masked[71];
  assign data_o[72] = data_masked[169] | data_masked[72];
  assign data_o[73] = data_masked[170] | data_masked[73];
  assign data_o[74] = data_masked[171] | data_masked[74];
  assign data_o[75] = data_masked[172] | data_masked[75];
  assign data_o[76] = data_masked[173] | data_masked[76];
  assign data_o[77] = data_masked[174] | data_masked[77];
  assign data_o[78] = data_masked[175] | data_masked[78];
  assign data_o[79] = data_masked[176] | data_masked[79];
  assign data_o[80] = data_masked[177] | data_masked[80];
  assign data_o[81] = data_masked[178] | data_masked[81];
  assign data_o[82] = data_masked[179] | data_masked[82];
  assign data_o[83] = data_masked[180] | data_masked[83];
  assign data_o[84] = data_masked[181] | data_masked[84];
  assign data_o[85] = data_masked[182] | data_masked[85];
  assign data_o[86] = data_masked[183] | data_masked[86];
  assign data_o[87] = data_masked[184] | data_masked[87];
  assign data_o[88] = data_masked[185] | data_masked[88];
  assign data_o[89] = data_masked[186] | data_masked[89];
  assign data_o[90] = data_masked[187] | data_masked[90];
  assign data_o[91] = data_masked[188] | data_masked[91];
  assign data_o[92] = data_masked[189] | data_masked[92];
  assign data_o[93] = data_masked[190] | data_masked[93];
  assign data_o[94] = data_masked[191] | data_masked[94];
  assign data_o[95] = data_masked[192] | data_masked[95];
  assign data_o[96] = data_masked[193] | data_masked[96];

endmodule



module bsg_unconcentrate_static_05_0
(
  i,
  o
);

  input [1:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_2_,o_0_;
  assign o[4] = 1'b0;
  assign o[3] = 1'b0;
  assign o[1] = 1'b0;
  assign o_2_ = i[1];
  assign o[2] = o_2_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_array_concentrate_static_03_97
(
  i,
  o
);

  input [484:0] i;
  output [193:0] o;
  wire [193:0] o;
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_03
(
  i,
  o
);

  input [4:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_unconcentrate_static_03_0
(
  i,
  o
);

  input [1:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_1_,o_0_;
  assign o[4] = 1'b0;
  assign o[3] = 1'b0;
  assign o[2] = 1'b0;
  assign o_1_ = i[1];
  assign o[1] = o_1_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_array_concentrate_static_17_97
(
  i,
  o
);

  input [484:0] i;
  output [387:0] o;
  wire [387:0] o;
  assign o[387] = i[484];
  assign o[386] = i[483];
  assign o[385] = i[482];
  assign o[384] = i[481];
  assign o[383] = i[480];
  assign o[382] = i[479];
  assign o[381] = i[478];
  assign o[380] = i[477];
  assign o[379] = i[476];
  assign o[378] = i[475];
  assign o[377] = i[474];
  assign o[376] = i[473];
  assign o[375] = i[472];
  assign o[374] = i[471];
  assign o[373] = i[470];
  assign o[372] = i[469];
  assign o[371] = i[468];
  assign o[370] = i[467];
  assign o[369] = i[466];
  assign o[368] = i[465];
  assign o[367] = i[464];
  assign o[366] = i[463];
  assign o[365] = i[462];
  assign o[364] = i[461];
  assign o[363] = i[460];
  assign o[362] = i[459];
  assign o[361] = i[458];
  assign o[360] = i[457];
  assign o[359] = i[456];
  assign o[358] = i[455];
  assign o[357] = i[454];
  assign o[356] = i[453];
  assign o[355] = i[452];
  assign o[354] = i[451];
  assign o[353] = i[450];
  assign o[352] = i[449];
  assign o[351] = i[448];
  assign o[350] = i[447];
  assign o[349] = i[446];
  assign o[348] = i[445];
  assign o[347] = i[444];
  assign o[346] = i[443];
  assign o[345] = i[442];
  assign o[344] = i[441];
  assign o[343] = i[440];
  assign o[342] = i[439];
  assign o[341] = i[438];
  assign o[340] = i[437];
  assign o[339] = i[436];
  assign o[338] = i[435];
  assign o[337] = i[434];
  assign o[336] = i[433];
  assign o[335] = i[432];
  assign o[334] = i[431];
  assign o[333] = i[430];
  assign o[332] = i[429];
  assign o[331] = i[428];
  assign o[330] = i[427];
  assign o[329] = i[426];
  assign o[328] = i[425];
  assign o[327] = i[424];
  assign o[326] = i[423];
  assign o[325] = i[422];
  assign o[324] = i[421];
  assign o[323] = i[420];
  assign o[322] = i[419];
  assign o[321] = i[418];
  assign o[320] = i[417];
  assign o[319] = i[416];
  assign o[318] = i[415];
  assign o[317] = i[414];
  assign o[316] = i[413];
  assign o[315] = i[412];
  assign o[314] = i[411];
  assign o[313] = i[410];
  assign o[312] = i[409];
  assign o[311] = i[408];
  assign o[310] = i[407];
  assign o[309] = i[406];
  assign o[308] = i[405];
  assign o[307] = i[404];
  assign o[306] = i[403];
  assign o[305] = i[402];
  assign o[304] = i[401];
  assign o[303] = i[400];
  assign o[302] = i[399];
  assign o[301] = i[398];
  assign o[300] = i[397];
  assign o[299] = i[396];
  assign o[298] = i[395];
  assign o[297] = i[394];
  assign o[296] = i[393];
  assign o[295] = i[392];
  assign o[294] = i[391];
  assign o[293] = i[390];
  assign o[292] = i[389];
  assign o[291] = i[388];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_17
(
  i,
  o
);

  input [4:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o[3] = i[4];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_scan_00000008_1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[7] | 1'b0;
  assign t_1__6_ = i[6] | i[7];
  assign t_1__5_ = i[5] | i[6];
  assign t_1__4_ = i[4] | i[5];
  assign t_1__3_ = i[3] | i[4];
  assign t_1__2_ = i[2] | i[3];
  assign t_1__1_ = i[1] | i[2];
  assign t_1__0_ = i[0] | i[1];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[7] = t_2__7_ | 1'b0;
  assign o[6] = t_2__6_ | 1'b0;
  assign o[5] = t_2__5_ | 1'b0;
  assign o[4] = t_2__4_ | 1'b0;
  assign o[3] = t_2__3_ | t_2__7_;
  assign o[2] = t_2__2_ | t_2__6_;
  assign o[1] = t_2__1_ | t_2__5_;
  assign o[0] = t_2__0_ | t_2__4_;

endmodule



module bsg_arb_round_robin_04
(
  clk_i,
  reset_i,
  reqs_i,
  grants_o,
  yumi_i
);

  input [3:0] reqs_i;
  output [3:0] grants_o;
  input clk_i;
  input reset_i;
  input yumi_i;
  wire [3:0] grants_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  wire [2:0] \fi2.thermocode_r ,\fi2.thermocode_n ;
  wire [6:4] \fi2.scan_li ;
  wire [7:0] \fi2.scan_lo ;
  wire [6:0] \fi2.edge_detect ;
  reg \fi2.thermocode_r_2_sv2v_reg ,\fi2.thermocode_r_1_sv2v_reg ,
  \fi2.thermocode_r_0_sv2v_reg ;
  assign \fi2.thermocode_r [2] = \fi2.thermocode_r_2_sv2v_reg ;
  assign \fi2.thermocode_r [1] = \fi2.thermocode_r_1_sv2v_reg ;
  assign \fi2.thermocode_r [0] = \fi2.thermocode_r_0_sv2v_reg ;

  bsg_scan_00000008_1
  \fi2.scan 
  (
    .i({ 1'b0, \fi2.scan_li , reqs_i }),
    .o(\fi2.scan_lo )
  );

  assign N3 = (N0)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = yumi_i;
  assign \fi2.thermocode_n  = (N1)? \fi2.scan_lo [7:5] : 
                              (N5)? \fi2.scan_lo [3:1] : 1'b0;
  assign N1 = N4;
  assign N2 = ~yumi_i;
  assign \fi2.scan_li [6] = \fi2.thermocode_r [2] & reqs_i[2];
  assign \fi2.scan_li [5] = \fi2.thermocode_r [1] & reqs_i[1];
  assign \fi2.scan_li [4] = \fi2.thermocode_r [0] & reqs_i[0];
  assign \fi2.edge_detect [6] = N6 & \fi2.scan_lo [6];
  assign N6 = ~\fi2.scan_lo [7];
  assign \fi2.edge_detect [5] = N7 & \fi2.scan_lo [5];
  assign N7 = ~\fi2.scan_lo [6];
  assign \fi2.edge_detect [4] = N8 & \fi2.scan_lo [4];
  assign N8 = ~\fi2.scan_lo [5];
  assign \fi2.edge_detect [3] = N9 & \fi2.scan_lo [3];
  assign N9 = ~\fi2.scan_lo [4];
  assign \fi2.edge_detect [2] = N10 & \fi2.scan_lo [2];
  assign N10 = ~\fi2.scan_lo [3];
  assign \fi2.edge_detect [1] = N11 & \fi2.scan_lo [1];
  assign N11 = ~\fi2.scan_lo [2];
  assign \fi2.edge_detect [0] = N12 & \fi2.scan_lo [0];
  assign N12 = ~\fi2.scan_lo [1];
  assign grants_o[3] = \fi2.scan_lo [7] | \fi2.edge_detect [3];
  assign grants_o[2] = \fi2.edge_detect [6] | \fi2.edge_detect [2];
  assign grants_o[1] = \fi2.edge_detect [5] | \fi2.edge_detect [1];
  assign grants_o[0] = \fi2.edge_detect [4] | \fi2.edge_detect [0];
  assign N4 = N14 | \fi2.scan_li [4];
  assign N14 = N13 | \fi2.scan_li [5];
  assign N13 = 1'b0 | \fi2.scan_li [6];
  assign N5 = ~N4;

  always @(posedge clk_i) begin
    if(reset_i) begin
      \fi2.thermocode_r_2_sv2v_reg  <= 1'b0;
      \fi2.thermocode_r_1_sv2v_reg  <= 1'b0;
      \fi2.thermocode_r_0_sv2v_reg  <= 1'b0;
    end else if(N3) begin
      \fi2.thermocode_r_2_sv2v_reg  <= \fi2.thermocode_n [2];
      \fi2.thermocode_r_1_sv2v_reg  <= \fi2.thermocode_n [1];
      \fi2.thermocode_r_0_sv2v_reg  <= \fi2.thermocode_n [0];
    end 
  end


endmodule



module bsg_mux_one_hot_97_04
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [387:0] data_i;
  input [3:0] sel_one_hot_i;
  output [96:0] data_o;
  wire [96:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193;
  wire [387:0] data_masked;
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[2];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[2];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[2];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[2];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[2];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[2];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[2];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[2];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[2];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[2];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[2];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[2];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[2];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[2];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[2];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[2];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[2];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[2];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[2];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[2];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[2];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[2];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[2];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[2];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[2];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[2];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[2];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[2];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[2];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[2];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[2];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[2];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[2];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[2];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[2];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[2];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[2];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[2];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[2];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[2];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[2];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[2];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[2];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[2];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[2];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[2];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[2];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[2];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[2];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[2];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[2];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[2];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[2];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[2];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[2];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[2];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[2];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[2];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[2];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[2];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[2];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[2];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[2];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[2];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[2];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[2];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[3];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[3];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[3];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[3];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[3];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[3];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[3];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[3];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[3];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[3];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[3];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[3];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[3];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[3];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[3];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[3];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[3];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[3];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[3];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[3];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[3];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[3];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[3];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[3];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[3];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[3];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[3];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[3];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[3];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[3];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[3];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[3];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[3];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[3];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[3];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[3];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[3];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[3];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[3];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[3];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[3];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[3];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[3];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[3];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[3];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[3];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[3];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[3];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[3];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[3];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[3];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[3];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[3];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[3];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[3];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[3];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[3];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[3];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[3];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[3];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[3];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[3];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[3];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[3];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[3];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[3];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[3];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[3];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[3];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[3];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[3];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[3];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[3];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[3];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[3];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[3];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[3];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[3];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[3];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[3];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[3];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[3];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[3];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[3];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[3];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[3];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[3];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[3];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[3];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[3];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[3];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[3];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[3];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[3];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[3];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[97];
  assign N0 = data_masked[291] | data_masked[194];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[98];
  assign N2 = data_masked[292] | data_masked[195];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[99];
  assign N4 = data_masked[293] | data_masked[196];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[100];
  assign N6 = data_masked[294] | data_masked[197];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[101];
  assign N8 = data_masked[295] | data_masked[198];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[102];
  assign N10 = data_masked[296] | data_masked[199];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[103];
  assign N12 = data_masked[297] | data_masked[200];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[104];
  assign N14 = data_masked[298] | data_masked[201];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[105];
  assign N16 = data_masked[299] | data_masked[202];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[106];
  assign N18 = data_masked[300] | data_masked[203];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[107];
  assign N20 = data_masked[301] | data_masked[204];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[108];
  assign N22 = data_masked[302] | data_masked[205];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[109];
  assign N24 = data_masked[303] | data_masked[206];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[110];
  assign N26 = data_masked[304] | data_masked[207];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[111];
  assign N28 = data_masked[305] | data_masked[208];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[112];
  assign N30 = data_masked[306] | data_masked[209];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[113];
  assign N32 = data_masked[307] | data_masked[210];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[114];
  assign N34 = data_masked[308] | data_masked[211];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[115];
  assign N36 = data_masked[309] | data_masked[212];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[116];
  assign N38 = data_masked[310] | data_masked[213];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[117];
  assign N40 = data_masked[311] | data_masked[214];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[118];
  assign N42 = data_masked[312] | data_masked[215];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[119];
  assign N44 = data_masked[313] | data_masked[216];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[120];
  assign N46 = data_masked[314] | data_masked[217];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[121];
  assign N48 = data_masked[315] | data_masked[218];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[122];
  assign N50 = data_masked[316] | data_masked[219];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[123];
  assign N52 = data_masked[317] | data_masked[220];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[124];
  assign N54 = data_masked[318] | data_masked[221];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[125];
  assign N56 = data_masked[319] | data_masked[222];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[126];
  assign N58 = data_masked[320] | data_masked[223];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[127];
  assign N60 = data_masked[321] | data_masked[224];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[128];
  assign N62 = data_masked[322] | data_masked[225];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[129];
  assign N64 = data_masked[323] | data_masked[226];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[130];
  assign N66 = data_masked[324] | data_masked[227];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[131];
  assign N68 = data_masked[325] | data_masked[228];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[132];
  assign N70 = data_masked[326] | data_masked[229];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[133];
  assign N72 = data_masked[327] | data_masked[230];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[134];
  assign N74 = data_masked[328] | data_masked[231];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[135];
  assign N76 = data_masked[329] | data_masked[232];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[136];
  assign N78 = data_masked[330] | data_masked[233];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[137];
  assign N80 = data_masked[331] | data_masked[234];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[138];
  assign N82 = data_masked[332] | data_masked[235];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[139];
  assign N84 = data_masked[333] | data_masked[236];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[140];
  assign N86 = data_masked[334] | data_masked[237];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[141];
  assign N88 = data_masked[335] | data_masked[238];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[142];
  assign N90 = data_masked[336] | data_masked[239];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[143];
  assign N92 = data_masked[337] | data_masked[240];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[144];
  assign N94 = data_masked[338] | data_masked[241];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[145];
  assign N96 = data_masked[339] | data_masked[242];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[146];
  assign N98 = data_masked[340] | data_masked[243];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[147];
  assign N100 = data_masked[341] | data_masked[244];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[148];
  assign N102 = data_masked[342] | data_masked[245];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[149];
  assign N104 = data_masked[343] | data_masked[246];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[150];
  assign N106 = data_masked[344] | data_masked[247];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[151];
  assign N108 = data_masked[345] | data_masked[248];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[152];
  assign N110 = data_masked[346] | data_masked[249];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[153];
  assign N112 = data_masked[347] | data_masked[250];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[154];
  assign N114 = data_masked[348] | data_masked[251];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[155];
  assign N116 = data_masked[349] | data_masked[252];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[156];
  assign N118 = data_masked[350] | data_masked[253];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[157];
  assign N120 = data_masked[351] | data_masked[254];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[158];
  assign N122 = data_masked[352] | data_masked[255];
  assign data_o[62] = N125 | data_masked[62];
  assign N125 = N124 | data_masked[159];
  assign N124 = data_masked[353] | data_masked[256];
  assign data_o[63] = N127 | data_masked[63];
  assign N127 = N126 | data_masked[160];
  assign N126 = data_masked[354] | data_masked[257];
  assign data_o[64] = N129 | data_masked[64];
  assign N129 = N128 | data_masked[161];
  assign N128 = data_masked[355] | data_masked[258];
  assign data_o[65] = N131 | data_masked[65];
  assign N131 = N130 | data_masked[162];
  assign N130 = data_masked[356] | data_masked[259];
  assign data_o[66] = N133 | data_masked[66];
  assign N133 = N132 | data_masked[163];
  assign N132 = data_masked[357] | data_masked[260];
  assign data_o[67] = N135 | data_masked[67];
  assign N135 = N134 | data_masked[164];
  assign N134 = data_masked[358] | data_masked[261];
  assign data_o[68] = N137 | data_masked[68];
  assign N137 = N136 | data_masked[165];
  assign N136 = data_masked[359] | data_masked[262];
  assign data_o[69] = N139 | data_masked[69];
  assign N139 = N138 | data_masked[166];
  assign N138 = data_masked[360] | data_masked[263];
  assign data_o[70] = N141 | data_masked[70];
  assign N141 = N140 | data_masked[167];
  assign N140 = data_masked[361] | data_masked[264];
  assign data_o[71] = N143 | data_masked[71];
  assign N143 = N142 | data_masked[168];
  assign N142 = data_masked[362] | data_masked[265];
  assign data_o[72] = N145 | data_masked[72];
  assign N145 = N144 | data_masked[169];
  assign N144 = data_masked[363] | data_masked[266];
  assign data_o[73] = N147 | data_masked[73];
  assign N147 = N146 | data_masked[170];
  assign N146 = data_masked[364] | data_masked[267];
  assign data_o[74] = N149 | data_masked[74];
  assign N149 = N148 | data_masked[171];
  assign N148 = data_masked[365] | data_masked[268];
  assign data_o[75] = N151 | data_masked[75];
  assign N151 = N150 | data_masked[172];
  assign N150 = data_masked[366] | data_masked[269];
  assign data_o[76] = N153 | data_masked[76];
  assign N153 = N152 | data_masked[173];
  assign N152 = data_masked[367] | data_masked[270];
  assign data_o[77] = N155 | data_masked[77];
  assign N155 = N154 | data_masked[174];
  assign N154 = data_masked[368] | data_masked[271];
  assign data_o[78] = N157 | data_masked[78];
  assign N157 = N156 | data_masked[175];
  assign N156 = data_masked[369] | data_masked[272];
  assign data_o[79] = N159 | data_masked[79];
  assign N159 = N158 | data_masked[176];
  assign N158 = data_masked[370] | data_masked[273];
  assign data_o[80] = N161 | data_masked[80];
  assign N161 = N160 | data_masked[177];
  assign N160 = data_masked[371] | data_masked[274];
  assign data_o[81] = N163 | data_masked[81];
  assign N163 = N162 | data_masked[178];
  assign N162 = data_masked[372] | data_masked[275];
  assign data_o[82] = N165 | data_masked[82];
  assign N165 = N164 | data_masked[179];
  assign N164 = data_masked[373] | data_masked[276];
  assign data_o[83] = N167 | data_masked[83];
  assign N167 = N166 | data_masked[180];
  assign N166 = data_masked[374] | data_masked[277];
  assign data_o[84] = N169 | data_masked[84];
  assign N169 = N168 | data_masked[181];
  assign N168 = data_masked[375] | data_masked[278];
  assign data_o[85] = N171 | data_masked[85];
  assign N171 = N170 | data_masked[182];
  assign N170 = data_masked[376] | data_masked[279];
  assign data_o[86] = N173 | data_masked[86];
  assign N173 = N172 | data_masked[183];
  assign N172 = data_masked[377] | data_masked[280];
  assign data_o[87] = N175 | data_masked[87];
  assign N175 = N174 | data_masked[184];
  assign N174 = data_masked[378] | data_masked[281];
  assign data_o[88] = N177 | data_masked[88];
  assign N177 = N176 | data_masked[185];
  assign N176 = data_masked[379] | data_masked[282];
  assign data_o[89] = N179 | data_masked[89];
  assign N179 = N178 | data_masked[186];
  assign N178 = data_masked[380] | data_masked[283];
  assign data_o[90] = N181 | data_masked[90];
  assign N181 = N180 | data_masked[187];
  assign N180 = data_masked[381] | data_masked[284];
  assign data_o[91] = N183 | data_masked[91];
  assign N183 = N182 | data_masked[188];
  assign N182 = data_masked[382] | data_masked[285];
  assign data_o[92] = N185 | data_masked[92];
  assign N185 = N184 | data_masked[189];
  assign N184 = data_masked[383] | data_masked[286];
  assign data_o[93] = N187 | data_masked[93];
  assign N187 = N186 | data_masked[190];
  assign N186 = data_masked[384] | data_masked[287];
  assign data_o[94] = N189 | data_masked[94];
  assign N189 = N188 | data_masked[191];
  assign N188 = data_masked[385] | data_masked[288];
  assign data_o[95] = N191 | data_masked[95];
  assign N191 = N190 | data_masked[192];
  assign N190 = data_masked[386] | data_masked[289];
  assign data_o[96] = N193 | data_masked[96];
  assign N193 = N192 | data_masked[193];
  assign N192 = data_masked[387] | data_masked[290];

endmodule



module bsg_unconcentrate_static_17_0
(
  i,
  o
);

  input [3:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_4_,o_2_,o_1_,o_0_;
  assign o[3] = 1'b0;
  assign o_4_ = i[3];
  assign o[4] = o_4_;
  assign o_2_ = i[2];
  assign o[2] = o_2_;
  assign o_1_ = i[1];
  assign o[1] = o_1_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_array_concentrate_static_0f_97
(
  i,
  o
);

  input [484:0] i;
  output [387:0] o;
  wire [387:0] o;
  assign o[387] = i[387];
  assign o[386] = i[386];
  assign o[385] = i[385];
  assign o[384] = i[384];
  assign o[383] = i[383];
  assign o[382] = i[382];
  assign o[381] = i[381];
  assign o[380] = i[380];
  assign o[379] = i[379];
  assign o[378] = i[378];
  assign o[377] = i[377];
  assign o[376] = i[376];
  assign o[375] = i[375];
  assign o[374] = i[374];
  assign o[373] = i[373];
  assign o[372] = i[372];
  assign o[371] = i[371];
  assign o[370] = i[370];
  assign o[369] = i[369];
  assign o[368] = i[368];
  assign o[367] = i[367];
  assign o[366] = i[366];
  assign o[365] = i[365];
  assign o[364] = i[364];
  assign o[363] = i[363];
  assign o[362] = i[362];
  assign o[361] = i[361];
  assign o[360] = i[360];
  assign o[359] = i[359];
  assign o[358] = i[358];
  assign o[357] = i[357];
  assign o[356] = i[356];
  assign o[355] = i[355];
  assign o[354] = i[354];
  assign o[353] = i[353];
  assign o[352] = i[352];
  assign o[351] = i[351];
  assign o[350] = i[350];
  assign o[349] = i[349];
  assign o[348] = i[348];
  assign o[347] = i[347];
  assign o[346] = i[346];
  assign o[345] = i[345];
  assign o[344] = i[344];
  assign o[343] = i[343];
  assign o[342] = i[342];
  assign o[341] = i[341];
  assign o[340] = i[340];
  assign o[339] = i[339];
  assign o[338] = i[338];
  assign o[337] = i[337];
  assign o[336] = i[336];
  assign o[335] = i[335];
  assign o[334] = i[334];
  assign o[333] = i[333];
  assign o[332] = i[332];
  assign o[331] = i[331];
  assign o[330] = i[330];
  assign o[329] = i[329];
  assign o[328] = i[328];
  assign o[327] = i[327];
  assign o[326] = i[326];
  assign o[325] = i[325];
  assign o[324] = i[324];
  assign o[323] = i[323];
  assign o[322] = i[322];
  assign o[321] = i[321];
  assign o[320] = i[320];
  assign o[319] = i[319];
  assign o[318] = i[318];
  assign o[317] = i[317];
  assign o[316] = i[316];
  assign o[315] = i[315];
  assign o[314] = i[314];
  assign o[313] = i[313];
  assign o[312] = i[312];
  assign o[311] = i[311];
  assign o[310] = i[310];
  assign o[309] = i[309];
  assign o[308] = i[308];
  assign o[307] = i[307];
  assign o[306] = i[306];
  assign o[305] = i[305];
  assign o[304] = i[304];
  assign o[303] = i[303];
  assign o[302] = i[302];
  assign o[301] = i[301];
  assign o[300] = i[300];
  assign o[299] = i[299];
  assign o[298] = i[298];
  assign o[297] = i[297];
  assign o[296] = i[296];
  assign o[295] = i[295];
  assign o[294] = i[294];
  assign o[293] = i[293];
  assign o[292] = i[292];
  assign o[291] = i[291];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_0f
(
  i,
  o
);

  input [4:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_unconcentrate_static_0f_0
(
  i,
  o
);

  input [3:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_3_,o_2_,o_1_,o_0_;
  assign o[4] = 1'b0;
  assign o_3_ = i[3];
  assign o[3] = o_3_;
  assign o_2_ = i[2];
  assign o[2] = o_2_;
  assign o_1_ = i[1];
  assign o[1] = o_1_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_mesh_router_width_p97_x_cord_width_p7_y_cord_width_p7_ruche_factor_X_p0_ruche_factor_Y_p0_dims_p2_XY_order_p1
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [484:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [484:0] data_o;
  output [4:0] v_o;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o,\dor_0_.temp_req ,\dor_1_.temp_req ,\dor_2_.temp_req ,
  \dor_3_.temp_req ,\dor_4_.temp_req ,\xbar_0_.conc_req ,\xbar_0_.grants ;
  wire [484:0] data_o,\xbar_0_.conc_data ;
  wire _0_net_,_1_net__4_,_1_net__3_,_1_net__2_,_1_net__1_,_1_net__0_,_2_net_,
  _3_net__1_,_3_net__0_,_4_net_,_5_net__1_,_5_net__0_,_6_net_,_7_net__3_,_7_net__2_,
  _7_net__1_,_7_net__0_,_8_net_,_9_net__3_,_9_net__2_,_9_net__1_,_9_net__0_,N0,N1,N2,N3,
  N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;
  wire [24:0] req,req_t,yumi_lo,yumi_lo_t;
  wire [193:0] \xbar_1_.conc_data ,\xbar_2_.conc_data ;
  wire [1:0] \xbar_1_.conc_req ,\xbar_1_.grants ,\xbar_2_.conc_req ,\xbar_2_.grants ;
  wire [387:0] \xbar_3_.conc_data ,\xbar_4_.conc_data ;
  wire [3:0] \xbar_3_.conc_req ,\xbar_3_.grants ,\xbar_4_.conc_req ,\xbar_4_.grants ;

  bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s01_0
  \dor_0_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[6:0]),
    .y_dirs_i(data_i[13:7]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_0_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s02_0
  \dor_1_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[103:97]),
    .y_dirs_i(data_i[110:104]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_1_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s04_0
  \dor_2_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[200:194]),
    .y_dirs_i(data_i[207:201]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_2_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s08_0
  \dor_3_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[297:291]),
    .y_dirs_i(data_i[304:298]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_3_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_1_s10_0
  \dor_4_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[394:388]),
    .y_dirs_i(data_i[401:395]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_4_.temp_req )
  );


  bsg_transpose_width_p5_els_p5
  req_tp
  (
    .i(req),
    .o(req_t)
  );


  bsg_array_concentrate_static_1f_97
  \xbar_0_.conc0 
  (
    .i(data_i),
    .o(\xbar_0_.conc_data )
  );


  bsg_concentrate_static_1f
  \xbar_0_.conc1 
  (
    .i(req_t[4:0]),
    .o(\xbar_0_.conc_req )
  );


  bsg_arb_round_robin_05
  \xbar_0_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_0_.conc_req ),
    .grants_o(\xbar_0_.grants ),
    .yumi_i(_0_net_)
  );


  bsg_mux_one_hot_97_05
  \xbar_0_.data_mux 
  (
    .data_i(\xbar_0_.conc_data ),
    .sel_one_hot_i(\xbar_0_.grants ),
    .data_o(data_o[96:0])
  );


  bsg_unconcentrate_static_1f_0
  \xbar_0_.unconc0 
  (
    .i({ _1_net__4_, _1_net__3_, _1_net__2_, _1_net__1_, _1_net__0_ }),
    .o(yumi_lo[4:0])
  );


  bsg_array_concentrate_static_05_97
  \xbar_1_.conc0 
  (
    .i(data_i),
    .o(\xbar_1_.conc_data )
  );


  bsg_concentrate_static_05
  \xbar_1_.conc1 
  (
    .i(req_t[9:5]),
    .o(\xbar_1_.conc_req )
  );


  bsg_arb_round_robin_02
  \xbar_1_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_1_.conc_req ),
    .grants_o(\xbar_1_.grants ),
    .yumi_i(_2_net_)
  );


  bsg_mux_one_hot_97_02
  \xbar_1_.data_mux 
  (
    .data_i(\xbar_1_.conc_data ),
    .sel_one_hot_i(\xbar_1_.grants ),
    .data_o(data_o[193:97])
  );


  bsg_unconcentrate_static_05_0
  \xbar_1_.unconc0 
  (
    .i({ _3_net__1_, _3_net__0_ }),
    .o(yumi_lo[9:5])
  );


  bsg_array_concentrate_static_03_97
  \xbar_2_.conc0 
  (
    .i(data_i),
    .o(\xbar_2_.conc_data )
  );


  bsg_concentrate_static_03
  \xbar_2_.conc1 
  (
    .i(req_t[14:10]),
    .o(\xbar_2_.conc_req )
  );


  bsg_arb_round_robin_02
  \xbar_2_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_2_.conc_req ),
    .grants_o(\xbar_2_.grants ),
    .yumi_i(_4_net_)
  );


  bsg_mux_one_hot_97_02
  \xbar_2_.data_mux 
  (
    .data_i(\xbar_2_.conc_data ),
    .sel_one_hot_i(\xbar_2_.grants ),
    .data_o(data_o[290:194])
  );


  bsg_unconcentrate_static_03_0
  \xbar_2_.unconc0 
  (
    .i({ _5_net__1_, _5_net__0_ }),
    .o(yumi_lo[14:10])
  );


  bsg_array_concentrate_static_17_97
  \xbar_3_.conc0 
  (
    .i(data_i),
    .o(\xbar_3_.conc_data )
  );


  bsg_concentrate_static_17
  \xbar_3_.conc1 
  (
    .i(req_t[19:15]),
    .o(\xbar_3_.conc_req )
  );


  bsg_arb_round_robin_04
  \xbar_3_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_3_.conc_req ),
    .grants_o(\xbar_3_.grants ),
    .yumi_i(_6_net_)
  );


  bsg_mux_one_hot_97_04
  \xbar_3_.data_mux 
  (
    .data_i(\xbar_3_.conc_data ),
    .sel_one_hot_i(\xbar_3_.grants ),
    .data_o(data_o[387:291])
  );


  bsg_unconcentrate_static_17_0
  \xbar_3_.unconc0 
  (
    .i({ _7_net__3_, _7_net__2_, _7_net__1_, _7_net__0_ }),
    .o(yumi_lo[19:15])
  );


  bsg_array_concentrate_static_0f_97
  \xbar_4_.conc0 
  (
    .i(data_i),
    .o(\xbar_4_.conc_data )
  );


  bsg_concentrate_static_0f
  \xbar_4_.conc1 
  (
    .i(req_t[24:20]),
    .o(\xbar_4_.conc_req )
  );


  bsg_arb_round_robin_04
  \xbar_4_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_4_.conc_req ),
    .grants_o(\xbar_4_.grants ),
    .yumi_i(_8_net_)
  );


  bsg_mux_one_hot_97_04
  \xbar_4_.data_mux 
  (
    .data_i(\xbar_4_.conc_data ),
    .sel_one_hot_i(\xbar_4_.grants ),
    .data_o(data_o[484:388])
  );


  bsg_unconcentrate_static_0f_0
  \xbar_4_.unconc0 
  (
    .i({ _9_net__3_, _9_net__2_, _9_net__1_, _9_net__0_ }),
    .o(yumi_lo[24:20])
  );


  bsg_transpose_width_p5_els_p5
  yumi_tp
  (
    .i(yumi_lo),
    .o(yumi_lo_t)
  );

  assign req[4] = v_i[0] & \dor_0_.temp_req [4];
  assign req[3] = v_i[0] & \dor_0_.temp_req [3];
  assign req[2] = v_i[0] & \dor_0_.temp_req [2];
  assign req[1] = v_i[0] & \dor_0_.temp_req [1];
  assign req[0] = v_i[0] & \dor_0_.temp_req [0];
  assign req[9] = v_i[1] & \dor_1_.temp_req [4];
  assign req[8] = v_i[1] & \dor_1_.temp_req [3];
  assign req[7] = v_i[1] & \dor_1_.temp_req [2];
  assign req[6] = v_i[1] & \dor_1_.temp_req [1];
  assign req[5] = v_i[1] & \dor_1_.temp_req [0];
  assign req[14] = v_i[2] & \dor_2_.temp_req [4];
  assign req[13] = v_i[2] & \dor_2_.temp_req [3];
  assign req[12] = v_i[2] & \dor_2_.temp_req [2];
  assign req[11] = v_i[2] & \dor_2_.temp_req [1];
  assign req[10] = v_i[2] & \dor_2_.temp_req [0];
  assign req[19] = v_i[3] & \dor_3_.temp_req [4];
  assign req[18] = v_i[3] & \dor_3_.temp_req [3];
  assign req[17] = v_i[3] & \dor_3_.temp_req [2];
  assign req[16] = v_i[3] & \dor_3_.temp_req [1];
  assign req[15] = v_i[3] & \dor_3_.temp_req [0];
  assign req[24] = v_i[4] & \dor_4_.temp_req [4];
  assign req[23] = v_i[4] & \dor_4_.temp_req [3];
  assign req[22] = v_i[4] & \dor_4_.temp_req [2];
  assign req[21] = v_i[4] & \dor_4_.temp_req [1];
  assign req[20] = v_i[4] & \dor_4_.temp_req [0];
  assign v_o[0] = N2 | \xbar_0_.conc_req [0];
  assign N2 = N1 | \xbar_0_.conc_req [1];
  assign N1 = N0 | \xbar_0_.conc_req [2];
  assign N0 = \xbar_0_.conc_req [4] | \xbar_0_.conc_req [3];
  assign _0_net_ = v_o[0] & ready_i[0];
  assign _1_net__4_ = \xbar_0_.grants [4] & ready_i[0];
  assign _1_net__3_ = \xbar_0_.grants [3] & ready_i[0];
  assign _1_net__2_ = \xbar_0_.grants [2] & ready_i[0];
  assign _1_net__1_ = \xbar_0_.grants [1] & ready_i[0];
  assign _1_net__0_ = \xbar_0_.grants [0] & ready_i[0];
  assign v_o[1] = \xbar_1_.conc_req [1] | \xbar_1_.conc_req [0];
  assign _2_net_ = v_o[1] & ready_i[1];
  assign _3_net__1_ = \xbar_1_.grants [1] & ready_i[1];
  assign _3_net__0_ = \xbar_1_.grants [0] & ready_i[1];
  assign v_o[2] = \xbar_2_.conc_req [1] | \xbar_2_.conc_req [0];
  assign _4_net_ = v_o[2] & ready_i[2];
  assign _5_net__1_ = \xbar_2_.grants [1] & ready_i[2];
  assign _5_net__0_ = \xbar_2_.grants [0] & ready_i[2];
  assign v_o[3] = N4 | \xbar_3_.conc_req [0];
  assign N4 = N3 | \xbar_3_.conc_req [1];
  assign N3 = \xbar_3_.conc_req [3] | \xbar_3_.conc_req [2];
  assign _6_net_ = v_o[3] & ready_i[3];
  assign _7_net__3_ = \xbar_3_.grants [3] & ready_i[3];
  assign _7_net__2_ = \xbar_3_.grants [2] & ready_i[3];
  assign _7_net__1_ = \xbar_3_.grants [1] & ready_i[3];
  assign _7_net__0_ = \xbar_3_.grants [0] & ready_i[3];
  assign v_o[4] = N6 | \xbar_4_.conc_req [0];
  assign N6 = N5 | \xbar_4_.conc_req [1];
  assign N5 = \xbar_4_.conc_req [3] | \xbar_4_.conc_req [2];
  assign _8_net_ = v_o[4] & ready_i[4];
  assign _9_net__3_ = \xbar_4_.grants [3] & ready_i[4];
  assign _9_net__2_ = \xbar_4_.grants [2] & ready_i[4];
  assign _9_net__1_ = \xbar_4_.grants [1] & ready_i[4];
  assign _9_net__0_ = \xbar_4_.grants [0] & ready_i[4];
  assign yumi_o[0] = N9 | yumi_lo_t[0];
  assign N9 = N8 | yumi_lo_t[1];
  assign N8 = N7 | yumi_lo_t[2];
  assign N7 = yumi_lo_t[4] | yumi_lo_t[3];
  assign yumi_o[1] = N12 | yumi_lo_t[5];
  assign N12 = N11 | yumi_lo_t[6];
  assign N11 = N10 | yumi_lo_t[7];
  assign N10 = yumi_lo_t[9] | yumi_lo_t[8];
  assign yumi_o[2] = N15 | yumi_lo_t[10];
  assign N15 = N14 | yumi_lo_t[11];
  assign N14 = N13 | yumi_lo_t[12];
  assign N13 = yumi_lo_t[14] | yumi_lo_t[13];
  assign yumi_o[3] = N18 | yumi_lo_t[15];
  assign N18 = N17 | yumi_lo_t[16];
  assign N17 = N16 | yumi_lo_t[17];
  assign N16 = yumi_lo_t[19] | yumi_lo_t[18];
  assign yumi_o[4] = N21 | yumi_lo_t[20];
  assign N21 = N20 | yumi_lo_t[21];
  assign N20 = N19 | yumi_lo_t[22];
  assign N19 = yumi_lo_t[24] | yumi_lo_t[23];

endmodule



module bsg_mesh_router_buffered_97_7_7_0_0_0_2_00_1_00_01
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [494:0] link_i;
  output [494:0] link_o;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [494:0] link_o;
  wire \rof_0_.fi.fifo_ready_lo ;
  wire [4:0] fifo_valid,fifo_yumi;
  wire [484:0] fifo_data;

  bsg_fifo_1r1w_small_width_p97_els_p3
  \rof_0_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[98]),
    .ready_o(\rof_0_.fi.fifo_ready_lo ),
    .data_i(link_i[96:0]),
    .v_o(fifo_valid[0]),
    .data_o(fifo_data[96:0]),
    .yumi_i(fifo_yumi[0])
  );


  bsg_dff_reset_width_p1_reset_val_p0
  \rof_0_.fi.cr.dff0 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(fifo_yumi[0]),
    .data_o(link_o[97])
  );


  bsg_fifo_1r1w_small_width_p97_els_p2
  \rof_1_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[197]),
    .ready_o(link_o[196]),
    .data_i(link_i[195:99]),
    .v_o(fifo_valid[1]),
    .data_o(fifo_data[193:97]),
    .yumi_i(fifo_yumi[1])
  );


  bsg_fifo_1r1w_small_width_p97_els_p2
  \rof_2_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[296]),
    .ready_o(link_o[295]),
    .data_i(link_i[294:198]),
    .v_o(fifo_valid[2]),
    .data_o(fifo_data[290:194]),
    .yumi_i(fifo_yumi[2])
  );


  bsg_fifo_1r1w_small_width_p97_els_p2
  \rof_3_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[395]),
    .ready_o(link_o[394]),
    .data_i(link_i[393:297]),
    .v_o(fifo_valid[3]),
    .data_o(fifo_data[387:291]),
    .yumi_i(fifo_yumi[3])
  );


  bsg_fifo_1r1w_small_width_p97_els_p2
  \rof_4_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[494]),
    .ready_o(link_o[493]),
    .data_i(link_i[492:396]),
    .v_o(fifo_valid[4]),
    .data_o(fifo_data[484:388]),
    .yumi_i(fifo_yumi[4])
  );


  bsg_mesh_router_width_p97_x_cord_width_p7_y_cord_width_p7_ruche_factor_X_p0_ruche_factor_Y_p0_dims_p2_XY_order_p1
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(fifo_data),
    .v_i(fifo_valid),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[493:493], link_i[394:394], link_i[295:295], link_i[196:196], link_i[97:97] }),
    .data_o({ link_o[492:396], link_o[393:297], link_o[294:198], link_o[195:99], link_o[96:0] }),
    .v_o({ link_o[494:494], link_o[395:395], link_o[296:296], link_o[197:197], link_o[98:98] }),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i)
  );


endmodule



module bsg_mem_1r1w_synth_width_p53_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [52:0] w_data_i;
  input [0:0] r_addr_i;
  output [52:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [52:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [105:0] \nz.mem ;
  reg \nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,
  \nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,
  \nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,
  \nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,
  \nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,
  \nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,
  \nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[52] = (N3)? \nz.mem [52] : 
                        (N0)? \nz.mem [105] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[51] = (N3)? \nz.mem [51] : 
                        (N0)? \nz.mem [104] : 1'b0;
  assign r_data_o[50] = (N3)? \nz.mem [50] : 
                        (N0)? \nz.mem [103] : 1'b0;
  assign r_data_o[49] = (N3)? \nz.mem [49] : 
                        (N0)? \nz.mem [102] : 1'b0;
  assign r_data_o[48] = (N3)? \nz.mem [48] : 
                        (N0)? \nz.mem [101] : 1'b0;
  assign r_data_o[47] = (N3)? \nz.mem [47] : 
                        (N0)? \nz.mem [100] : 1'b0;
  assign r_data_o[46] = (N3)? \nz.mem [46] : 
                        (N0)? \nz.mem [99] : 1'b0;
  assign r_data_o[45] = (N3)? \nz.mem [45] : 
                        (N0)? \nz.mem [98] : 1'b0;
  assign r_data_o[44] = (N3)? \nz.mem [44] : 
                        (N0)? \nz.mem [97] : 1'b0;
  assign r_data_o[43] = (N3)? \nz.mem [43] : 
                        (N0)? \nz.mem [96] : 1'b0;
  assign r_data_o[42] = (N3)? \nz.mem [42] : 
                        (N0)? \nz.mem [95] : 1'b0;
  assign r_data_o[41] = (N3)? \nz.mem [41] : 
                        (N0)? \nz.mem [94] : 1'b0;
  assign r_data_o[40] = (N3)? \nz.mem [40] : 
                        (N0)? \nz.mem [93] : 1'b0;
  assign r_data_o[39] = (N3)? \nz.mem [39] : 
                        (N0)? \nz.mem [92] : 1'b0;
  assign r_data_o[38] = (N3)? \nz.mem [38] : 
                        (N0)? \nz.mem [91] : 1'b0;
  assign r_data_o[37] = (N3)? \nz.mem [37] : 
                        (N0)? \nz.mem [90] : 1'b0;
  assign r_data_o[36] = (N3)? \nz.mem [36] : 
                        (N0)? \nz.mem [89] : 1'b0;
  assign r_data_o[35] = (N3)? \nz.mem [35] : 
                        (N0)? \nz.mem [88] : 1'b0;
  assign r_data_o[34] = (N3)? \nz.mem [34] : 
                        (N0)? \nz.mem [87] : 1'b0;
  assign r_data_o[33] = (N3)? \nz.mem [33] : 
                        (N0)? \nz.mem [86] : 1'b0;
  assign r_data_o[32] = (N3)? \nz.mem [32] : 
                        (N0)? \nz.mem [85] : 1'b0;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [84] : 1'b0;
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [83] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [82] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [81] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [80] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [79] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [78] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [77] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [76] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [75] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [74] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [73] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [72] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [71] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [70] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [69] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [68] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [67] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [66] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [65] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [64] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [63] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [62] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [61] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [60] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [59] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [58] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [57] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [56] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [55] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [54] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [53] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_105_sv2v_reg  <= w_data_i[52];
      \nz.mem_104_sv2v_reg  <= w_data_i[51];
      \nz.mem_103_sv2v_reg  <= w_data_i[50];
      \nz.mem_102_sv2v_reg  <= w_data_i[49];
      \nz.mem_101_sv2v_reg  <= w_data_i[48];
      \nz.mem_100_sv2v_reg  <= w_data_i[47];
      \nz.mem_99_sv2v_reg  <= w_data_i[46];
      \nz.mem_98_sv2v_reg  <= w_data_i[45];
      \nz.mem_97_sv2v_reg  <= w_data_i[44];
      \nz.mem_96_sv2v_reg  <= w_data_i[43];
      \nz.mem_95_sv2v_reg  <= w_data_i[42];
      \nz.mem_94_sv2v_reg  <= w_data_i[41];
      \nz.mem_93_sv2v_reg  <= w_data_i[40];
      \nz.mem_92_sv2v_reg  <= w_data_i[39];
      \nz.mem_91_sv2v_reg  <= w_data_i[38];
      \nz.mem_90_sv2v_reg  <= w_data_i[37];
      \nz.mem_89_sv2v_reg  <= w_data_i[36];
      \nz.mem_88_sv2v_reg  <= w_data_i[35];
      \nz.mem_87_sv2v_reg  <= w_data_i[34];
      \nz.mem_86_sv2v_reg  <= w_data_i[33];
      \nz.mem_85_sv2v_reg  <= w_data_i[32];
      \nz.mem_84_sv2v_reg  <= w_data_i[31];
      \nz.mem_83_sv2v_reg  <= w_data_i[30];
      \nz.mem_82_sv2v_reg  <= w_data_i[29];
      \nz.mem_81_sv2v_reg  <= w_data_i[28];
      \nz.mem_80_sv2v_reg  <= w_data_i[27];
      \nz.mem_79_sv2v_reg  <= w_data_i[26];
      \nz.mem_78_sv2v_reg  <= w_data_i[25];
      \nz.mem_77_sv2v_reg  <= w_data_i[24];
      \nz.mem_76_sv2v_reg  <= w_data_i[23];
      \nz.mem_75_sv2v_reg  <= w_data_i[22];
      \nz.mem_74_sv2v_reg  <= w_data_i[21];
      \nz.mem_73_sv2v_reg  <= w_data_i[20];
      \nz.mem_72_sv2v_reg  <= w_data_i[19];
      \nz.mem_71_sv2v_reg  <= w_data_i[18];
      \nz.mem_70_sv2v_reg  <= w_data_i[17];
      \nz.mem_69_sv2v_reg  <= w_data_i[16];
      \nz.mem_68_sv2v_reg  <= w_data_i[15];
      \nz.mem_67_sv2v_reg  <= w_data_i[14];
      \nz.mem_66_sv2v_reg  <= w_data_i[13];
      \nz.mem_65_sv2v_reg  <= w_data_i[12];
      \nz.mem_64_sv2v_reg  <= w_data_i[11];
      \nz.mem_63_sv2v_reg  <= w_data_i[10];
      \nz.mem_62_sv2v_reg  <= w_data_i[9];
      \nz.mem_61_sv2v_reg  <= w_data_i[8];
      \nz.mem_60_sv2v_reg  <= w_data_i[7];
      \nz.mem_59_sv2v_reg  <= w_data_i[6];
      \nz.mem_58_sv2v_reg  <= w_data_i[5];
      \nz.mem_57_sv2v_reg  <= w_data_i[4];
      \nz.mem_56_sv2v_reg  <= w_data_i[3];
      \nz.mem_55_sv2v_reg  <= w_data_i[2];
      \nz.mem_54_sv2v_reg  <= w_data_i[1];
      \nz.mem_53_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p53_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [52:0] w_data_i;
  input [0:0] r_addr_i;
  output [52:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [52:0] r_data_o;

  bsg_mem_1r1w_synth_width_p53_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p53_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [52:0] data_i;
  output [52:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [52:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p53_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_fifo_1r1w_small_width_p53_els_p2
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [52:0] data_i;
  output [52:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [52:0] data_o;
  wire ready_o,v_o;

  bsg_two_fifo_width_p53_ready_THEN_valid_p0
  \unhardened.tf.twof 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_i(v_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s01_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,x_gt,x_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign x_gt = x_dirs_i > my_x_i;
  assign req_o[4] = y_dirs_i > my_y_i;
  assign x_lt = N0 & N1;
  assign N0 = ~x_gt;
  assign N1 = ~x_eq;
  assign req_o[3] = N2 & N3;
  assign N2 = ~req_o[4];
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[1] = y_eq & x_lt;
  assign req_o[2] = y_eq & x_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s02_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,x_gt,x_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign x_gt = x_dirs_i > my_x_i;
  assign req_o[4] = y_dirs_i > my_y_i;
  assign x_lt = N0 & N1;
  assign N0 = ~x_gt;
  assign N1 = ~x_eq;
  assign req_o[3] = N2 & N3;
  assign N2 = ~req_o[4];
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[1] = y_eq & x_lt;
  assign req_o[2] = y_eq & x_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s04_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,x_gt,x_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign x_gt = x_dirs_i > my_x_i;
  assign req_o[4] = y_dirs_i > my_y_i;
  assign x_lt = N0 & N1;
  assign N0 = ~x_gt;
  assign N1 = ~x_eq;
  assign req_o[3] = N2 & N3;
  assign N2 = ~req_o[4];
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[1] = y_eq & x_lt;
  assign req_o[2] = y_eq & x_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s08_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,x_gt,x_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign x_gt = x_dirs_i > my_x_i;
  assign req_o[4] = y_dirs_i > my_y_i;
  assign x_lt = N0 & N1;
  assign N0 = ~x_gt;
  assign N1 = ~x_eq;
  assign req_o[3] = N2 & N3;
  assign N2 = ~req_o[4];
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[1] = y_eq & x_lt;
  assign req_o[2] = y_eq & x_gt;

endmodule



module bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s10_0
(
  clk_i,
  reset_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [6:0] x_dirs_i;
  input [6:0] y_dirs_i;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  output [4:0] req_o;
  input clk_i;
  input reset_i;
  wire [4:0] req_o;
  wire x_eq,y_eq,x_gt,x_lt,N0,N1,N2,N3;
  assign x_eq = x_dirs_i == my_x_i;
  assign y_eq = y_dirs_i == my_y_i;
  assign x_gt = x_dirs_i > my_x_i;
  assign req_o[4] = y_dirs_i > my_y_i;
  assign x_lt = N0 & N1;
  assign N0 = ~x_gt;
  assign N1 = ~x_eq;
  assign req_o[3] = N2 & N3;
  assign N2 = ~req_o[4];
  assign N3 = ~y_eq;
  assign req_o[0] = x_eq & y_eq;
  assign req_o[1] = y_eq & x_lt;
  assign req_o[2] = y_eq & x_gt;

endmodule



module bsg_array_concentrate_static_1f_53
(
  i,
  o
);

  input [264:0] i;
  output [264:0] o;
  wire [264:0] o;
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_mux_one_hot_53_05
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [264:0] data_i;
  input [4:0] sel_one_hot_i;
  output [52:0] data_o;
  wire [52:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158;
  wire [264:0] data_masked;
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[2];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[2];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[2];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[2];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[2];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[2];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[2];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[2];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[2];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[2];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[2];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[2];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[2];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[2];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[2];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[2];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[2];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[2];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[2];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[2];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[2];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[3];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[3];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[3];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[3];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[3];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[3];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[3];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[3];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[3];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[3];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[3];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[3];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[3];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[3];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[3];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[3];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[3];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[3];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[3];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[3];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[3];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[3];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[3];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[3];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[3];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[3];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[3];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[3];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[3];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[3];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[3];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[3];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[3];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[4];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[4];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[4];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[4];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[4];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[4];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[4];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[4];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[4];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[4];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[4];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[4];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[4];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[4];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[4];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[4];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[4];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[4];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[4];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[4];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[4];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[4];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[4];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[4];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[4];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[4];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[4];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[4];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[4];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[4];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[4];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[4];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[4];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[4];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[4];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[4];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[4];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[4];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[4];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[4];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[4];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[4];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[4];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[53];
  assign N1 = N0 | data_masked[106];
  assign N0 = data_masked[212] | data_masked[159];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[54];
  assign N4 = N3 | data_masked[107];
  assign N3 = data_masked[213] | data_masked[160];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[55];
  assign N7 = N6 | data_masked[108];
  assign N6 = data_masked[214] | data_masked[161];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[56];
  assign N10 = N9 | data_masked[109];
  assign N9 = data_masked[215] | data_masked[162];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[57];
  assign N13 = N12 | data_masked[110];
  assign N12 = data_masked[216] | data_masked[163];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[58];
  assign N16 = N15 | data_masked[111];
  assign N15 = data_masked[217] | data_masked[164];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[59];
  assign N19 = N18 | data_masked[112];
  assign N18 = data_masked[218] | data_masked[165];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[60];
  assign N22 = N21 | data_masked[113];
  assign N21 = data_masked[219] | data_masked[166];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[61];
  assign N25 = N24 | data_masked[114];
  assign N24 = data_masked[220] | data_masked[167];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[62];
  assign N28 = N27 | data_masked[115];
  assign N27 = data_masked[221] | data_masked[168];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[63];
  assign N31 = N30 | data_masked[116];
  assign N30 = data_masked[222] | data_masked[169];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[64];
  assign N34 = N33 | data_masked[117];
  assign N33 = data_masked[223] | data_masked[170];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[65];
  assign N37 = N36 | data_masked[118];
  assign N36 = data_masked[224] | data_masked[171];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[66];
  assign N40 = N39 | data_masked[119];
  assign N39 = data_masked[225] | data_masked[172];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[67];
  assign N43 = N42 | data_masked[120];
  assign N42 = data_masked[226] | data_masked[173];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[68];
  assign N46 = N45 | data_masked[121];
  assign N45 = data_masked[227] | data_masked[174];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[69];
  assign N49 = N48 | data_masked[122];
  assign N48 = data_masked[228] | data_masked[175];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[70];
  assign N52 = N51 | data_masked[123];
  assign N51 = data_masked[229] | data_masked[176];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[71];
  assign N55 = N54 | data_masked[124];
  assign N54 = data_masked[230] | data_masked[177];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[72];
  assign N58 = N57 | data_masked[125];
  assign N57 = data_masked[231] | data_masked[178];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[73];
  assign N61 = N60 | data_masked[126];
  assign N60 = data_masked[232] | data_masked[179];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[74];
  assign N64 = N63 | data_masked[127];
  assign N63 = data_masked[233] | data_masked[180];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[75];
  assign N67 = N66 | data_masked[128];
  assign N66 = data_masked[234] | data_masked[181];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[76];
  assign N70 = N69 | data_masked[129];
  assign N69 = data_masked[235] | data_masked[182];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[77];
  assign N73 = N72 | data_masked[130];
  assign N72 = data_masked[236] | data_masked[183];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[78];
  assign N76 = N75 | data_masked[131];
  assign N75 = data_masked[237] | data_masked[184];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[79];
  assign N79 = N78 | data_masked[132];
  assign N78 = data_masked[238] | data_masked[185];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[80];
  assign N82 = N81 | data_masked[133];
  assign N81 = data_masked[239] | data_masked[186];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[81];
  assign N85 = N84 | data_masked[134];
  assign N84 = data_masked[240] | data_masked[187];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[82];
  assign N88 = N87 | data_masked[135];
  assign N87 = data_masked[241] | data_masked[188];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[83];
  assign N91 = N90 | data_masked[136];
  assign N90 = data_masked[242] | data_masked[189];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[84];
  assign N94 = N93 | data_masked[137];
  assign N93 = data_masked[243] | data_masked[190];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[85];
  assign N97 = N96 | data_masked[138];
  assign N96 = data_masked[244] | data_masked[191];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[86];
  assign N100 = N99 | data_masked[139];
  assign N99 = data_masked[245] | data_masked[192];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[87];
  assign N103 = N102 | data_masked[140];
  assign N102 = data_masked[246] | data_masked[193];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[88];
  assign N106 = N105 | data_masked[141];
  assign N105 = data_masked[247] | data_masked[194];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[89];
  assign N109 = N108 | data_masked[142];
  assign N108 = data_masked[248] | data_masked[195];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[90];
  assign N112 = N111 | data_masked[143];
  assign N111 = data_masked[249] | data_masked[196];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[91];
  assign N115 = N114 | data_masked[144];
  assign N114 = data_masked[250] | data_masked[197];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[92];
  assign N118 = N117 | data_masked[145];
  assign N117 = data_masked[251] | data_masked[198];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[93];
  assign N121 = N120 | data_masked[146];
  assign N120 = data_masked[252] | data_masked[199];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[94];
  assign N124 = N123 | data_masked[147];
  assign N123 = data_masked[253] | data_masked[200];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[95];
  assign N127 = N126 | data_masked[148];
  assign N126 = data_masked[254] | data_masked[201];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[96];
  assign N130 = N129 | data_masked[149];
  assign N129 = data_masked[255] | data_masked[202];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[97];
  assign N133 = N132 | data_masked[150];
  assign N132 = data_masked[256] | data_masked[203];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[98];
  assign N136 = N135 | data_masked[151];
  assign N135 = data_masked[257] | data_masked[204];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[99];
  assign N139 = N138 | data_masked[152];
  assign N138 = data_masked[258] | data_masked[205];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[100];
  assign N142 = N141 | data_masked[153];
  assign N141 = data_masked[259] | data_masked[206];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[101];
  assign N145 = N144 | data_masked[154];
  assign N144 = data_masked[260] | data_masked[207];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[102];
  assign N148 = N147 | data_masked[155];
  assign N147 = data_masked[261] | data_masked[208];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[103];
  assign N151 = N150 | data_masked[156];
  assign N150 = data_masked[262] | data_masked[209];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[104];
  assign N154 = N153 | data_masked[157];
  assign N153 = data_masked[263] | data_masked[210];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[105];
  assign N157 = N156 | data_masked[158];
  assign N156 = data_masked[264] | data_masked[211];

endmodule



module bsg_array_concentrate_static_1d_53
(
  i,
  o
);

  input [264:0] i;
  output [211:0] o;
  wire [211:0] o;
  assign o[211] = i[264];
  assign o[210] = i[263];
  assign o[209] = i[262];
  assign o[208] = i[261];
  assign o[207] = i[260];
  assign o[206] = i[259];
  assign o[205] = i[258];
  assign o[204] = i[257];
  assign o[203] = i[256];
  assign o[202] = i[255];
  assign o[201] = i[254];
  assign o[200] = i[253];
  assign o[199] = i[252];
  assign o[198] = i[251];
  assign o[197] = i[250];
  assign o[196] = i[249];
  assign o[195] = i[248];
  assign o[194] = i[247];
  assign o[193] = i[246];
  assign o[192] = i[245];
  assign o[191] = i[244];
  assign o[190] = i[243];
  assign o[189] = i[242];
  assign o[188] = i[241];
  assign o[187] = i[240];
  assign o[186] = i[239];
  assign o[185] = i[238];
  assign o[184] = i[237];
  assign o[183] = i[236];
  assign o[182] = i[235];
  assign o[181] = i[234];
  assign o[180] = i[233];
  assign o[179] = i[232];
  assign o[178] = i[231];
  assign o[177] = i[230];
  assign o[176] = i[229];
  assign o[175] = i[228];
  assign o[174] = i[227];
  assign o[173] = i[226];
  assign o[172] = i[225];
  assign o[171] = i[224];
  assign o[170] = i[223];
  assign o[169] = i[222];
  assign o[168] = i[221];
  assign o[167] = i[220];
  assign o[166] = i[219];
  assign o[165] = i[218];
  assign o[164] = i[217];
  assign o[163] = i[216];
  assign o[162] = i[215];
  assign o[161] = i[214];
  assign o[160] = i[213];
  assign o[159] = i[212];
  assign o[158] = i[211];
  assign o[157] = i[210];
  assign o[156] = i[209];
  assign o[155] = i[208];
  assign o[154] = i[207];
  assign o[153] = i[206];
  assign o[152] = i[205];
  assign o[151] = i[204];
  assign o[150] = i[203];
  assign o[149] = i[202];
  assign o[148] = i[201];
  assign o[147] = i[200];
  assign o[146] = i[199];
  assign o[145] = i[198];
  assign o[144] = i[197];
  assign o[143] = i[196];
  assign o[142] = i[195];
  assign o[141] = i[194];
  assign o[140] = i[193];
  assign o[139] = i[192];
  assign o[138] = i[191];
  assign o[137] = i[190];
  assign o[136] = i[189];
  assign o[135] = i[188];
  assign o[134] = i[187];
  assign o[133] = i[186];
  assign o[132] = i[185];
  assign o[131] = i[184];
  assign o[130] = i[183];
  assign o[129] = i[182];
  assign o[128] = i[181];
  assign o[127] = i[180];
  assign o[126] = i[179];
  assign o[125] = i[178];
  assign o[124] = i[177];
  assign o[123] = i[176];
  assign o[122] = i[175];
  assign o[121] = i[174];
  assign o[120] = i[173];
  assign o[119] = i[172];
  assign o[118] = i[171];
  assign o[117] = i[170];
  assign o[116] = i[169];
  assign o[115] = i[168];
  assign o[114] = i[167];
  assign o[113] = i[166];
  assign o[112] = i[165];
  assign o[111] = i[164];
  assign o[110] = i[163];
  assign o[109] = i[162];
  assign o[108] = i[161];
  assign o[107] = i[160];
  assign o[106] = i[159];
  assign o[105] = i[158];
  assign o[104] = i[157];
  assign o[103] = i[156];
  assign o[102] = i[155];
  assign o[101] = i[154];
  assign o[100] = i[153];
  assign o[99] = i[152];
  assign o[98] = i[151];
  assign o[97] = i[150];
  assign o[96] = i[149];
  assign o[95] = i[148];
  assign o[94] = i[147];
  assign o[93] = i[146];
  assign o[92] = i[145];
  assign o[91] = i[144];
  assign o[90] = i[143];
  assign o[89] = i[142];
  assign o[88] = i[141];
  assign o[87] = i[140];
  assign o[86] = i[139];
  assign o[85] = i[138];
  assign o[84] = i[137];
  assign o[83] = i[136];
  assign o[82] = i[135];
  assign o[81] = i[134];
  assign o[80] = i[133];
  assign o[79] = i[132];
  assign o[78] = i[131];
  assign o[77] = i[130];
  assign o[76] = i[129];
  assign o[75] = i[128];
  assign o[74] = i[127];
  assign o[73] = i[126];
  assign o[72] = i[125];
  assign o[71] = i[124];
  assign o[70] = i[123];
  assign o[69] = i[122];
  assign o[68] = i[121];
  assign o[67] = i[120];
  assign o[66] = i[119];
  assign o[65] = i[118];
  assign o[64] = i[117];
  assign o[63] = i[116];
  assign o[62] = i[115];
  assign o[61] = i[114];
  assign o[60] = i[113];
  assign o[59] = i[112];
  assign o[58] = i[111];
  assign o[57] = i[110];
  assign o[56] = i[109];
  assign o[55] = i[108];
  assign o[54] = i[107];
  assign o[53] = i[106];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_1d
(
  i,
  o
);

  input [4:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o[3] = i[4];
  assign o[2] = i[3];
  assign o[1] = i[2];
  assign o[0] = i[0];

endmodule



module bsg_mux_one_hot_53_04
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [211:0] data_i;
  input [3:0] sel_one_hot_i;
  output [52:0] data_o;
  wire [52:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105;
  wire [211:0] data_masked;
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[2];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[2];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[2];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[2];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[2];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[2];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[2];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[2];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[2];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[2];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[2];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[2];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[2];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[2];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[2];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[2];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[2];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[2];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[2];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[2];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[2];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[3];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[3];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[3];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[3];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[3];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[3];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[3];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[3];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[3];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[3];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[3];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[3];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[3];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[3];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[3];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[3];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[3];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[3];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[3];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[3];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[3];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[3];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[3];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[3];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[3];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[3];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[3];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[3];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[3];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[3];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[3];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[3];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[53];
  assign N0 = data_masked[159] | data_masked[106];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[54];
  assign N2 = data_masked[160] | data_masked[107];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[55];
  assign N4 = data_masked[161] | data_masked[108];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[56];
  assign N6 = data_masked[162] | data_masked[109];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[57];
  assign N8 = data_masked[163] | data_masked[110];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[58];
  assign N10 = data_masked[164] | data_masked[111];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[59];
  assign N12 = data_masked[165] | data_masked[112];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[60];
  assign N14 = data_masked[166] | data_masked[113];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[61];
  assign N16 = data_masked[167] | data_masked[114];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[62];
  assign N18 = data_masked[168] | data_masked[115];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[63];
  assign N20 = data_masked[169] | data_masked[116];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[64];
  assign N22 = data_masked[170] | data_masked[117];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[65];
  assign N24 = data_masked[171] | data_masked[118];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[66];
  assign N26 = data_masked[172] | data_masked[119];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[67];
  assign N28 = data_masked[173] | data_masked[120];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[68];
  assign N30 = data_masked[174] | data_masked[121];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[69];
  assign N32 = data_masked[175] | data_masked[122];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[70];
  assign N34 = data_masked[176] | data_masked[123];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[71];
  assign N36 = data_masked[177] | data_masked[124];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[72];
  assign N38 = data_masked[178] | data_masked[125];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[73];
  assign N40 = data_masked[179] | data_masked[126];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[74];
  assign N42 = data_masked[180] | data_masked[127];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[75];
  assign N44 = data_masked[181] | data_masked[128];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[76];
  assign N46 = data_masked[182] | data_masked[129];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[77];
  assign N48 = data_masked[183] | data_masked[130];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[78];
  assign N50 = data_masked[184] | data_masked[131];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[79];
  assign N52 = data_masked[185] | data_masked[132];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[80];
  assign N54 = data_masked[186] | data_masked[133];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[81];
  assign N56 = data_masked[187] | data_masked[134];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[82];
  assign N58 = data_masked[188] | data_masked[135];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[83];
  assign N60 = data_masked[189] | data_masked[136];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[84];
  assign N62 = data_masked[190] | data_masked[137];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[85];
  assign N64 = data_masked[191] | data_masked[138];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[86];
  assign N66 = data_masked[192] | data_masked[139];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[87];
  assign N68 = data_masked[193] | data_masked[140];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[88];
  assign N70 = data_masked[194] | data_masked[141];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[89];
  assign N72 = data_masked[195] | data_masked[142];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[90];
  assign N74 = data_masked[196] | data_masked[143];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[91];
  assign N76 = data_masked[197] | data_masked[144];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[92];
  assign N78 = data_masked[198] | data_masked[145];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[93];
  assign N80 = data_masked[199] | data_masked[146];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[94];
  assign N82 = data_masked[200] | data_masked[147];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[95];
  assign N84 = data_masked[201] | data_masked[148];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[96];
  assign N86 = data_masked[202] | data_masked[149];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[97];
  assign N88 = data_masked[203] | data_masked[150];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[98];
  assign N90 = data_masked[204] | data_masked[151];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[99];
  assign N92 = data_masked[205] | data_masked[152];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[100];
  assign N94 = data_masked[206] | data_masked[153];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[101];
  assign N96 = data_masked[207] | data_masked[154];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[102];
  assign N98 = data_masked[208] | data_masked[155];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[103];
  assign N100 = data_masked[209] | data_masked[156];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[104];
  assign N102 = data_masked[210] | data_masked[157];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[105];
  assign N104 = data_masked[211] | data_masked[158];

endmodule



module bsg_unconcentrate_static_1d_0
(
  i,
  o
);

  input [3:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_4_,o_3_,o_2_,o_0_;
  assign o[1] = 1'b0;
  assign o_4_ = i[3];
  assign o[4] = o_4_;
  assign o_3_ = i[2];
  assign o[3] = o_3_;
  assign o_2_ = i[1];
  assign o[2] = o_2_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_array_concentrate_static_1b_53
(
  i,
  o
);

  input [264:0] i;
  output [211:0] o;
  wire [211:0] o;
  assign o[211] = i[264];
  assign o[210] = i[263];
  assign o[209] = i[262];
  assign o[208] = i[261];
  assign o[207] = i[260];
  assign o[206] = i[259];
  assign o[205] = i[258];
  assign o[204] = i[257];
  assign o[203] = i[256];
  assign o[202] = i[255];
  assign o[201] = i[254];
  assign o[200] = i[253];
  assign o[199] = i[252];
  assign o[198] = i[251];
  assign o[197] = i[250];
  assign o[196] = i[249];
  assign o[195] = i[248];
  assign o[194] = i[247];
  assign o[193] = i[246];
  assign o[192] = i[245];
  assign o[191] = i[244];
  assign o[190] = i[243];
  assign o[189] = i[242];
  assign o[188] = i[241];
  assign o[187] = i[240];
  assign o[186] = i[239];
  assign o[185] = i[238];
  assign o[184] = i[237];
  assign o[183] = i[236];
  assign o[182] = i[235];
  assign o[181] = i[234];
  assign o[180] = i[233];
  assign o[179] = i[232];
  assign o[178] = i[231];
  assign o[177] = i[230];
  assign o[176] = i[229];
  assign o[175] = i[228];
  assign o[174] = i[227];
  assign o[173] = i[226];
  assign o[172] = i[225];
  assign o[171] = i[224];
  assign o[170] = i[223];
  assign o[169] = i[222];
  assign o[168] = i[221];
  assign o[167] = i[220];
  assign o[166] = i[219];
  assign o[165] = i[218];
  assign o[164] = i[217];
  assign o[163] = i[216];
  assign o[162] = i[215];
  assign o[161] = i[214];
  assign o[160] = i[213];
  assign o[159] = i[212];
  assign o[158] = i[211];
  assign o[157] = i[210];
  assign o[156] = i[209];
  assign o[155] = i[208];
  assign o[154] = i[207];
  assign o[153] = i[206];
  assign o[152] = i[205];
  assign o[151] = i[204];
  assign o[150] = i[203];
  assign o[149] = i[202];
  assign o[148] = i[201];
  assign o[147] = i[200];
  assign o[146] = i[199];
  assign o[145] = i[198];
  assign o[144] = i[197];
  assign o[143] = i[196];
  assign o[142] = i[195];
  assign o[141] = i[194];
  assign o[140] = i[193];
  assign o[139] = i[192];
  assign o[138] = i[191];
  assign o[137] = i[190];
  assign o[136] = i[189];
  assign o[135] = i[188];
  assign o[134] = i[187];
  assign o[133] = i[186];
  assign o[132] = i[185];
  assign o[131] = i[184];
  assign o[130] = i[183];
  assign o[129] = i[182];
  assign o[128] = i[181];
  assign o[127] = i[180];
  assign o[126] = i[179];
  assign o[125] = i[178];
  assign o[124] = i[177];
  assign o[123] = i[176];
  assign o[122] = i[175];
  assign o[121] = i[174];
  assign o[120] = i[173];
  assign o[119] = i[172];
  assign o[118] = i[171];
  assign o[117] = i[170];
  assign o[116] = i[169];
  assign o[115] = i[168];
  assign o[114] = i[167];
  assign o[113] = i[166];
  assign o[112] = i[165];
  assign o[111] = i[164];
  assign o[110] = i[163];
  assign o[109] = i[162];
  assign o[108] = i[161];
  assign o[107] = i[160];
  assign o[106] = i[159];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_1b
(
  i,
  o
);

  input [4:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o[3] = i[4];
  assign o[2] = i[3];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_unconcentrate_static_1b_0
(
  i,
  o
);

  input [3:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_4_,o_3_,o_1_,o_0_;
  assign o[2] = 1'b0;
  assign o_4_ = i[3];
  assign o[4] = o_4_;
  assign o_3_ = i[2];
  assign o[3] = o_3_;
  assign o_1_ = i[1];
  assign o[1] = o_1_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_array_concentrate_static_11_53
(
  i,
  o
);

  input [264:0] i;
  output [105:0] o;
  wire [105:0] o;
  assign o[105] = i[264];
  assign o[104] = i[263];
  assign o[103] = i[262];
  assign o[102] = i[261];
  assign o[101] = i[260];
  assign o[100] = i[259];
  assign o[99] = i[258];
  assign o[98] = i[257];
  assign o[97] = i[256];
  assign o[96] = i[255];
  assign o[95] = i[254];
  assign o[94] = i[253];
  assign o[93] = i[252];
  assign o[92] = i[251];
  assign o[91] = i[250];
  assign o[90] = i[249];
  assign o[89] = i[248];
  assign o[88] = i[247];
  assign o[87] = i[246];
  assign o[86] = i[245];
  assign o[85] = i[244];
  assign o[84] = i[243];
  assign o[83] = i[242];
  assign o[82] = i[241];
  assign o[81] = i[240];
  assign o[80] = i[239];
  assign o[79] = i[238];
  assign o[78] = i[237];
  assign o[77] = i[236];
  assign o[76] = i[235];
  assign o[75] = i[234];
  assign o[74] = i[233];
  assign o[73] = i[232];
  assign o[72] = i[231];
  assign o[71] = i[230];
  assign o[70] = i[229];
  assign o[69] = i[228];
  assign o[68] = i[227];
  assign o[67] = i[226];
  assign o[66] = i[225];
  assign o[65] = i[224];
  assign o[64] = i[223];
  assign o[63] = i[222];
  assign o[62] = i[221];
  assign o[61] = i[220];
  assign o[60] = i[219];
  assign o[59] = i[218];
  assign o[58] = i[217];
  assign o[57] = i[216];
  assign o[56] = i[215];
  assign o[55] = i[214];
  assign o[54] = i[213];
  assign o[53] = i[212];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_11
(
  i,
  o
);

  input [4:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[1] = i[4];
  assign o[0] = i[0];

endmodule



module bsg_mux_one_hot_53_02
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [105:0] data_i;
  input [1:0] sel_one_hot_i;
  output [52:0] data_o;
  wire [52:0] data_o;
  wire [105:0] data_masked;
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[53] | data_masked[0];
  assign data_o[1] = data_masked[54] | data_masked[1];
  assign data_o[2] = data_masked[55] | data_masked[2];
  assign data_o[3] = data_masked[56] | data_masked[3];
  assign data_o[4] = data_masked[57] | data_masked[4];
  assign data_o[5] = data_masked[58] | data_masked[5];
  assign data_o[6] = data_masked[59] | data_masked[6];
  assign data_o[7] = data_masked[60] | data_masked[7];
  assign data_o[8] = data_masked[61] | data_masked[8];
  assign data_o[9] = data_masked[62] | data_masked[9];
  assign data_o[10] = data_masked[63] | data_masked[10];
  assign data_o[11] = data_masked[64] | data_masked[11];
  assign data_o[12] = data_masked[65] | data_masked[12];
  assign data_o[13] = data_masked[66] | data_masked[13];
  assign data_o[14] = data_masked[67] | data_masked[14];
  assign data_o[15] = data_masked[68] | data_masked[15];
  assign data_o[16] = data_masked[69] | data_masked[16];
  assign data_o[17] = data_masked[70] | data_masked[17];
  assign data_o[18] = data_masked[71] | data_masked[18];
  assign data_o[19] = data_masked[72] | data_masked[19];
  assign data_o[20] = data_masked[73] | data_masked[20];
  assign data_o[21] = data_masked[74] | data_masked[21];
  assign data_o[22] = data_masked[75] | data_masked[22];
  assign data_o[23] = data_masked[76] | data_masked[23];
  assign data_o[24] = data_masked[77] | data_masked[24];
  assign data_o[25] = data_masked[78] | data_masked[25];
  assign data_o[26] = data_masked[79] | data_masked[26];
  assign data_o[27] = data_masked[80] | data_masked[27];
  assign data_o[28] = data_masked[81] | data_masked[28];
  assign data_o[29] = data_masked[82] | data_masked[29];
  assign data_o[30] = data_masked[83] | data_masked[30];
  assign data_o[31] = data_masked[84] | data_masked[31];
  assign data_o[32] = data_masked[85] | data_masked[32];
  assign data_o[33] = data_masked[86] | data_masked[33];
  assign data_o[34] = data_masked[87] | data_masked[34];
  assign data_o[35] = data_masked[88] | data_masked[35];
  assign data_o[36] = data_masked[89] | data_masked[36];
  assign data_o[37] = data_masked[90] | data_masked[37];
  assign data_o[38] = data_masked[91] | data_masked[38];
  assign data_o[39] = data_masked[92] | data_masked[39];
  assign data_o[40] = data_masked[93] | data_masked[40];
  assign data_o[41] = data_masked[94] | data_masked[41];
  assign data_o[42] = data_masked[95] | data_masked[42];
  assign data_o[43] = data_masked[96] | data_masked[43];
  assign data_o[44] = data_masked[97] | data_masked[44];
  assign data_o[45] = data_masked[98] | data_masked[45];
  assign data_o[46] = data_masked[99] | data_masked[46];
  assign data_o[47] = data_masked[100] | data_masked[47];
  assign data_o[48] = data_masked[101] | data_masked[48];
  assign data_o[49] = data_masked[102] | data_masked[49];
  assign data_o[50] = data_masked[103] | data_masked[50];
  assign data_o[51] = data_masked[104] | data_masked[51];
  assign data_o[52] = data_masked[105] | data_masked[52];

endmodule



module bsg_unconcentrate_static_11_0
(
  i,
  o
);

  input [1:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_4_,o_0_;
  assign o[3] = 1'b0;
  assign o[2] = 1'b0;
  assign o[1] = 1'b0;
  assign o_4_ = i[1];
  assign o[4] = o_4_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_array_concentrate_static_09_53
(
  i,
  o
);

  input [264:0] i;
  output [105:0] o;
  wire [105:0] o;
  assign o[105] = i[211];
  assign o[104] = i[210];
  assign o[103] = i[209];
  assign o[102] = i[208];
  assign o[101] = i[207];
  assign o[100] = i[206];
  assign o[99] = i[205];
  assign o[98] = i[204];
  assign o[97] = i[203];
  assign o[96] = i[202];
  assign o[95] = i[201];
  assign o[94] = i[200];
  assign o[93] = i[199];
  assign o[92] = i[198];
  assign o[91] = i[197];
  assign o[90] = i[196];
  assign o[89] = i[195];
  assign o[88] = i[194];
  assign o[87] = i[193];
  assign o[86] = i[192];
  assign o[85] = i[191];
  assign o[84] = i[190];
  assign o[83] = i[189];
  assign o[82] = i[188];
  assign o[81] = i[187];
  assign o[80] = i[186];
  assign o[79] = i[185];
  assign o[78] = i[184];
  assign o[77] = i[183];
  assign o[76] = i[182];
  assign o[75] = i[181];
  assign o[74] = i[180];
  assign o[73] = i[179];
  assign o[72] = i[178];
  assign o[71] = i[177];
  assign o[70] = i[176];
  assign o[69] = i[175];
  assign o[68] = i[174];
  assign o[67] = i[173];
  assign o[66] = i[172];
  assign o[65] = i[171];
  assign o[64] = i[170];
  assign o[63] = i[169];
  assign o[62] = i[168];
  assign o[61] = i[167];
  assign o[60] = i[166];
  assign o[59] = i[165];
  assign o[58] = i[164];
  assign o[57] = i[163];
  assign o[56] = i[162];
  assign o[55] = i[161];
  assign o[54] = i[160];
  assign o[53] = i[159];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_concentrate_static_09
(
  i,
  o
);

  input [4:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[1] = i[3];
  assign o[0] = i[0];

endmodule



module bsg_unconcentrate_static_09_0
(
  i,
  o
);

  input [1:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire o_3_,o_0_;
  assign o[4] = 1'b0;
  assign o[2] = 1'b0;
  assign o[1] = 1'b0;
  assign o_3_ = i[1];
  assign o[3] = o_3_;
  assign o_0_ = i[0];
  assign o[0] = o_0_;

endmodule



module bsg_mesh_router_width_p53_x_cord_width_p7_y_cord_width_p7_ruche_factor_X_p0_ruche_factor_Y_p0_dims_p2_XY_order_p0
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [264:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [264:0] data_o;
  output [4:0] v_o;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o,\dor_0_.temp_req ,\dor_1_.temp_req ,\dor_2_.temp_req ,
  \dor_3_.temp_req ,\dor_4_.temp_req ,\xbar_0_.conc_req ,\xbar_0_.grants ;
  wire [264:0] data_o,\xbar_0_.conc_data ;
  wire _0_net_,_1_net__4_,_1_net__3_,_1_net__2_,_1_net__1_,_1_net__0_,_2_net_,
  _3_net__3_,_3_net__2_,_3_net__1_,_3_net__0_,_4_net_,_5_net__3_,_5_net__2_,_5_net__1_,
  _5_net__0_,_6_net_,_7_net__1_,_7_net__0_,_8_net_,_9_net__1_,_9_net__0_,N0,N1,N2,N3,
  N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;
  wire [24:0] req,req_t,yumi_lo,yumi_lo_t;
  wire [211:0] \xbar_1_.conc_data ,\xbar_2_.conc_data ;
  wire [3:0] \xbar_1_.conc_req ,\xbar_1_.grants ,\xbar_2_.conc_req ,\xbar_2_.grants ;
  wire [105:0] \xbar_3_.conc_data ,\xbar_4_.conc_data ;
  wire [1:0] \xbar_3_.conc_req ,\xbar_3_.grants ,\xbar_4_.conc_req ,\xbar_4_.grants ;

  bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s01_0
  \dor_0_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[6:0]),
    .y_dirs_i(data_i[13:7]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_0_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s02_0
  \dor_1_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[59:53]),
    .y_dirs_i(data_i[66:60]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_1_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s04_0
  \dor_2_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[112:106]),
    .y_dirs_i(data_i[119:113]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_2_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s08_0
  \dor_3_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[165:159]),
    .y_dirs_i(data_i[172:166]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_3_.temp_req )
  );


  bsg_mesh_router_decoder_dor_7_7_2_0_0_0_s10_0
  \dor_4_.dor_decoder 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .x_dirs_i(data_i[218:212]),
    .y_dirs_i(data_i[225:219]),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .req_o(\dor_4_.temp_req )
  );


  bsg_transpose_width_p5_els_p5
  req_tp
  (
    .i(req),
    .o(req_t)
  );


  bsg_array_concentrate_static_1f_53
  \xbar_0_.conc0 
  (
    .i(data_i),
    .o(\xbar_0_.conc_data )
  );


  bsg_concentrate_static_1f
  \xbar_0_.conc1 
  (
    .i(req_t[4:0]),
    .o(\xbar_0_.conc_req )
  );


  bsg_arb_round_robin_05
  \xbar_0_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_0_.conc_req ),
    .grants_o(\xbar_0_.grants ),
    .yumi_i(_0_net_)
  );


  bsg_mux_one_hot_53_05
  \xbar_0_.data_mux 
  (
    .data_i(\xbar_0_.conc_data ),
    .sel_one_hot_i(\xbar_0_.grants ),
    .data_o(data_o[52:0])
  );


  bsg_unconcentrate_static_1f_0
  \xbar_0_.unconc0 
  (
    .i({ _1_net__4_, _1_net__3_, _1_net__2_, _1_net__1_, _1_net__0_ }),
    .o(yumi_lo[4:0])
  );


  bsg_array_concentrate_static_1d_53
  \xbar_1_.conc0 
  (
    .i(data_i),
    .o(\xbar_1_.conc_data )
  );


  bsg_concentrate_static_1d
  \xbar_1_.conc1 
  (
    .i(req_t[9:5]),
    .o(\xbar_1_.conc_req )
  );


  bsg_arb_round_robin_04
  \xbar_1_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_1_.conc_req ),
    .grants_o(\xbar_1_.grants ),
    .yumi_i(_2_net_)
  );


  bsg_mux_one_hot_53_04
  \xbar_1_.data_mux 
  (
    .data_i(\xbar_1_.conc_data ),
    .sel_one_hot_i(\xbar_1_.grants ),
    .data_o(data_o[105:53])
  );


  bsg_unconcentrate_static_1d_0
  \xbar_1_.unconc0 
  (
    .i({ _3_net__3_, _3_net__2_, _3_net__1_, _3_net__0_ }),
    .o(yumi_lo[9:5])
  );


  bsg_array_concentrate_static_1b_53
  \xbar_2_.conc0 
  (
    .i(data_i),
    .o(\xbar_2_.conc_data )
  );


  bsg_concentrate_static_1b
  \xbar_2_.conc1 
  (
    .i(req_t[14:10]),
    .o(\xbar_2_.conc_req )
  );


  bsg_arb_round_robin_04
  \xbar_2_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_2_.conc_req ),
    .grants_o(\xbar_2_.grants ),
    .yumi_i(_4_net_)
  );


  bsg_mux_one_hot_53_04
  \xbar_2_.data_mux 
  (
    .data_i(\xbar_2_.conc_data ),
    .sel_one_hot_i(\xbar_2_.grants ),
    .data_o(data_o[158:106])
  );


  bsg_unconcentrate_static_1b_0
  \xbar_2_.unconc0 
  (
    .i({ _5_net__3_, _5_net__2_, _5_net__1_, _5_net__0_ }),
    .o(yumi_lo[14:10])
  );


  bsg_array_concentrate_static_11_53
  \xbar_3_.conc0 
  (
    .i(data_i),
    .o(\xbar_3_.conc_data )
  );


  bsg_concentrate_static_11
  \xbar_3_.conc1 
  (
    .i(req_t[19:15]),
    .o(\xbar_3_.conc_req )
  );


  bsg_arb_round_robin_02
  \xbar_3_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_3_.conc_req ),
    .grants_o(\xbar_3_.grants ),
    .yumi_i(_6_net_)
  );


  bsg_mux_one_hot_53_02
  \xbar_3_.data_mux 
  (
    .data_i(\xbar_3_.conc_data ),
    .sel_one_hot_i(\xbar_3_.grants ),
    .data_o(data_o[211:159])
  );


  bsg_unconcentrate_static_11_0
  \xbar_3_.unconc0 
  (
    .i({ _7_net__1_, _7_net__0_ }),
    .o(yumi_lo[19:15])
  );


  bsg_array_concentrate_static_09_53
  \xbar_4_.conc0 
  (
    .i(data_i),
    .o(\xbar_4_.conc_data )
  );


  bsg_concentrate_static_09
  \xbar_4_.conc1 
  (
    .i(req_t[24:20]),
    .o(\xbar_4_.conc_req )
  );


  bsg_arb_round_robin_02
  \xbar_4_.rr 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .reqs_i(\xbar_4_.conc_req ),
    .grants_o(\xbar_4_.grants ),
    .yumi_i(_8_net_)
  );


  bsg_mux_one_hot_53_02
  \xbar_4_.data_mux 
  (
    .data_i(\xbar_4_.conc_data ),
    .sel_one_hot_i(\xbar_4_.grants ),
    .data_o(data_o[264:212])
  );


  bsg_unconcentrate_static_09_0
  \xbar_4_.unconc0 
  (
    .i({ _9_net__1_, _9_net__0_ }),
    .o(yumi_lo[24:20])
  );


  bsg_transpose_width_p5_els_p5
  yumi_tp
  (
    .i(yumi_lo),
    .o(yumi_lo_t)
  );

  assign req[4] = v_i[0] & \dor_0_.temp_req [4];
  assign req[3] = v_i[0] & \dor_0_.temp_req [3];
  assign req[2] = v_i[0] & \dor_0_.temp_req [2];
  assign req[1] = v_i[0] & \dor_0_.temp_req [1];
  assign req[0] = v_i[0] & \dor_0_.temp_req [0];
  assign req[9] = v_i[1] & \dor_1_.temp_req [4];
  assign req[8] = v_i[1] & \dor_1_.temp_req [3];
  assign req[7] = v_i[1] & \dor_1_.temp_req [2];
  assign req[6] = v_i[1] & \dor_1_.temp_req [1];
  assign req[5] = v_i[1] & \dor_1_.temp_req [0];
  assign req[14] = v_i[2] & \dor_2_.temp_req [4];
  assign req[13] = v_i[2] & \dor_2_.temp_req [3];
  assign req[12] = v_i[2] & \dor_2_.temp_req [2];
  assign req[11] = v_i[2] & \dor_2_.temp_req [1];
  assign req[10] = v_i[2] & \dor_2_.temp_req [0];
  assign req[19] = v_i[3] & \dor_3_.temp_req [4];
  assign req[18] = v_i[3] & \dor_3_.temp_req [3];
  assign req[17] = v_i[3] & \dor_3_.temp_req [2];
  assign req[16] = v_i[3] & \dor_3_.temp_req [1];
  assign req[15] = v_i[3] & \dor_3_.temp_req [0];
  assign req[24] = v_i[4] & \dor_4_.temp_req [4];
  assign req[23] = v_i[4] & \dor_4_.temp_req [3];
  assign req[22] = v_i[4] & \dor_4_.temp_req [2];
  assign req[21] = v_i[4] & \dor_4_.temp_req [1];
  assign req[20] = v_i[4] & \dor_4_.temp_req [0];
  assign v_o[0] = N2 | \xbar_0_.conc_req [0];
  assign N2 = N1 | \xbar_0_.conc_req [1];
  assign N1 = N0 | \xbar_0_.conc_req [2];
  assign N0 = \xbar_0_.conc_req [4] | \xbar_0_.conc_req [3];
  assign _0_net_ = v_o[0] & ready_i[0];
  assign _1_net__4_ = \xbar_0_.grants [4] & ready_i[0];
  assign _1_net__3_ = \xbar_0_.grants [3] & ready_i[0];
  assign _1_net__2_ = \xbar_0_.grants [2] & ready_i[0];
  assign _1_net__1_ = \xbar_0_.grants [1] & ready_i[0];
  assign _1_net__0_ = \xbar_0_.grants [0] & ready_i[0];
  assign v_o[1] = N4 | \xbar_1_.conc_req [0];
  assign N4 = N3 | \xbar_1_.conc_req [1];
  assign N3 = \xbar_1_.conc_req [3] | \xbar_1_.conc_req [2];
  assign _2_net_ = v_o[1] & ready_i[1];
  assign _3_net__3_ = \xbar_1_.grants [3] & ready_i[1];
  assign _3_net__2_ = \xbar_1_.grants [2] & ready_i[1];
  assign _3_net__1_ = \xbar_1_.grants [1] & ready_i[1];
  assign _3_net__0_ = \xbar_1_.grants [0] & ready_i[1];
  assign v_o[2] = N6 | \xbar_2_.conc_req [0];
  assign N6 = N5 | \xbar_2_.conc_req [1];
  assign N5 = \xbar_2_.conc_req [3] | \xbar_2_.conc_req [2];
  assign _4_net_ = v_o[2] & ready_i[2];
  assign _5_net__3_ = \xbar_2_.grants [3] & ready_i[2];
  assign _5_net__2_ = \xbar_2_.grants [2] & ready_i[2];
  assign _5_net__1_ = \xbar_2_.grants [1] & ready_i[2];
  assign _5_net__0_ = \xbar_2_.grants [0] & ready_i[2];
  assign v_o[3] = \xbar_3_.conc_req [1] | \xbar_3_.conc_req [0];
  assign _6_net_ = v_o[3] & ready_i[3];
  assign _7_net__1_ = \xbar_3_.grants [1] & ready_i[3];
  assign _7_net__0_ = \xbar_3_.grants [0] & ready_i[3];
  assign v_o[4] = \xbar_4_.conc_req [1] | \xbar_4_.conc_req [0];
  assign _8_net_ = v_o[4] & ready_i[4];
  assign _9_net__1_ = \xbar_4_.grants [1] & ready_i[4];
  assign _9_net__0_ = \xbar_4_.grants [0] & ready_i[4];
  assign yumi_o[0] = N9 | yumi_lo_t[0];
  assign N9 = N8 | yumi_lo_t[1];
  assign N8 = N7 | yumi_lo_t[2];
  assign N7 = yumi_lo_t[4] | yumi_lo_t[3];
  assign yumi_o[1] = N12 | yumi_lo_t[5];
  assign N12 = N11 | yumi_lo_t[6];
  assign N11 = N10 | yumi_lo_t[7];
  assign N10 = yumi_lo_t[9] | yumi_lo_t[8];
  assign yumi_o[2] = N15 | yumi_lo_t[10];
  assign N15 = N14 | yumi_lo_t[11];
  assign N14 = N13 | yumi_lo_t[12];
  assign N13 = yumi_lo_t[14] | yumi_lo_t[13];
  assign yumi_o[3] = N18 | yumi_lo_t[15];
  assign N18 = N17 | yumi_lo_t[16];
  assign N17 = N16 | yumi_lo_t[17];
  assign N16 = yumi_lo_t[19] | yumi_lo_t[18];
  assign yumi_o[4] = N21 | yumi_lo_t[20];
  assign N21 = N20 | yumi_lo_t[21];
  assign N20 = N19 | yumi_lo_t[22];
  assign N19 = yumi_lo_t[24] | yumi_lo_t[23];

endmodule



module bsg_mesh_router_buffered_53_7_7_0_0_0_2_00_0_00_00
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [274:0] link_i;
  output [274:0] link_o;
  input [6:0] my_x_i;
  input [6:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [274:0] link_o;
  wire [4:0] fifo_valid,fifo_yumi;
  wire [264:0] fifo_data;

  bsg_fifo_1r1w_small_width_p53_els_p2
  \rof_0_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[54]),
    .ready_o(link_o[53]),
    .data_i(link_i[52:0]),
    .v_o(fifo_valid[0]),
    .data_o(fifo_data[52:0]),
    .yumi_i(fifo_yumi[0])
  );


  bsg_fifo_1r1w_small_width_p53_els_p2
  \rof_1_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[109]),
    .ready_o(link_o[108]),
    .data_i(link_i[107:55]),
    .v_o(fifo_valid[1]),
    .data_o(fifo_data[105:53]),
    .yumi_i(fifo_yumi[1])
  );


  bsg_fifo_1r1w_small_width_p53_els_p2
  \rof_2_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[164]),
    .ready_o(link_o[163]),
    .data_i(link_i[162:110]),
    .v_o(fifo_valid[2]),
    .data_o(fifo_data[158:106]),
    .yumi_i(fifo_yumi[2])
  );


  bsg_fifo_1r1w_small_width_p53_els_p2
  \rof_3_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[219]),
    .ready_o(link_o[218]),
    .data_i(link_i[217:165]),
    .v_o(fifo_valid[3]),
    .data_o(fifo_data[211:159]),
    .yumi_i(fifo_yumi[3])
  );


  bsg_fifo_1r1w_small_width_p53_els_p2
  \rof_4_.fi.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_i[274]),
    .ready_o(link_o[273]),
    .data_i(link_i[272:220]),
    .v_o(fifo_valid[4]),
    .data_o(fifo_data[264:212]),
    .yumi_i(fifo_yumi[4])
  );


  bsg_mesh_router_width_p53_x_cord_width_p7_y_cord_width_p7_ruche_factor_X_p0_ruche_factor_Y_p0_dims_p2_XY_order_p0
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(fifo_data),
    .v_i(fifo_valid),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[273:273], link_i[218:218], link_i[163:163], link_i[108:108], link_i[53:53] }),
    .data_o({ link_o[272:220], link_o[217:165], link_o[162:110], link_o[107:55], link_o[52:0] }),
    .v_o({ link_o[274:274], link_o[219:219], link_o[164:164], link_o[109:109], link_o[54:54] }),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i)
  );


endmodule



module bsg_manycore_mesh_node_7_7_32_28_2_0_0_01_00_0
(
  clk_i,
  reset_i,
  links_sif_i,
  links_sif_o,
  proc_link_sif_i,
  proc_link_sif_o,
  global_x_i,
  global_y_i
);

  input [615:0] links_sif_i;
  output [615:0] links_sif_o;
  input [153:0] proc_link_sif_i;
  output [153:0] proc_link_sif_o;
  input [6:0] global_x_i;
  input [6:0] global_y_i;
  input clk_i;
  input reset_i;
  wire [615:0] links_sif_o;
  wire [153:0] proc_link_sif_o;

  bsg_mesh_router_buffered_97_7_7_0_0_0_2_00_1_00_01
  fwd
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ links_sif_i[615:517], links_sif_i[461:363], links_sif_i[307:209], links_sif_i[153:55], proc_link_sif_i[153:55] }),
    .link_o({ links_sif_o[615:517], links_sif_o[461:363], links_sif_o[307:209], links_sif_o[153:55], proc_link_sif_o[153:55] }),
    .my_x_i(global_x_i),
    .my_y_i(global_y_i)
  );


  bsg_mesh_router_buffered_53_7_7_0_0_0_2_00_0_00_00
  rev
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ links_sif_i[516:462], links_sif_i[362:308], links_sif_i[208:154], links_sif_i[54:0], proc_link_sif_i[54:0] }),
    .link_o({ links_sif_o[516:462], links_sif_o[362:308], links_sif_o[208:154], links_sif_o[54:0], proc_link_sif_o[54:0] }),
    .my_x_i(global_x_i),
    .my_y_i(global_y_i)
  );


endmodule



module bsg_circular_ptr_slots_p4_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1  = o + 1'b1;
  assign n_o = (N0)? \genblk1.genblk1.ptr_r_p1  : 
               (N1)? o : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_els_p4
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,N0,N1,N2,enq_r,deq_r,N3,equal_ptrs,sv2v_dc_1,sv2v_dc_2;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_slots_p4_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p4_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N3 = (N0)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = N1;
  assign N1 = enq_i | deq_i;
  assign N2 = ~N1;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N3) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p97_els_p4_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [96:0] w_data_i;
  input [1:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;
  wire [387:0] \nz.mem ;
  reg \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,
  \nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,
  \nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,
  \nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,
  \nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,
  \nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,
  \nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,
  \nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,
  \nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,
  \nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,
  \nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,
  \nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,
  \nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,
  \nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,
  \nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,
  \nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,
  \nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,
  \nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,
  \nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,
  \nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,
  \nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,
  \nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,
  \nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,
  \nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,
  \nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,
  \nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,
  \nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,
  \nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,
  \nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,
  \nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,
  \nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,
  \nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,
  \nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,
  \nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,
  \nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,
  \nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,
  \nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,
  \nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,
  \nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,
  \nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,
  \nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,
  \nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,
  \nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,
  \nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,
  \nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,
  \nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,
  \nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,
  \nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,
  \nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,
  \nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,
  \nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,
  \nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,
  \nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,
  \nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,
  \nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,
  \nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,
  \nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,
  \nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,
  \nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,
  \nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,
  \nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,
  \nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,
  \nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,
  \nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,
  \nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,
  \nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,
  \nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,
  \nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,
  \nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,
  \nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,
  \nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,
  \nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,
  \nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,
  \nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[96] = (N8)? \nz.mem [96] : 
                        (N10)? \nz.mem [193] : 
                        (N9)? \nz.mem [290] : 
                        (N11)? \nz.mem [387] : 1'b0;
  assign r_data_o[95] = (N8)? \nz.mem [95] : 
                        (N10)? \nz.mem [192] : 
                        (N9)? \nz.mem [289] : 
                        (N11)? \nz.mem [386] : 1'b0;
  assign r_data_o[94] = (N8)? \nz.mem [94] : 
                        (N10)? \nz.mem [191] : 
                        (N9)? \nz.mem [288] : 
                        (N11)? \nz.mem [385] : 1'b0;
  assign r_data_o[93] = (N8)? \nz.mem [93] : 
                        (N10)? \nz.mem [190] : 
                        (N9)? \nz.mem [287] : 
                        (N11)? \nz.mem [384] : 1'b0;
  assign r_data_o[92] = (N8)? \nz.mem [92] : 
                        (N10)? \nz.mem [189] : 
                        (N9)? \nz.mem [286] : 
                        (N11)? \nz.mem [383] : 1'b0;
  assign r_data_o[91] = (N8)? \nz.mem [91] : 
                        (N10)? \nz.mem [188] : 
                        (N9)? \nz.mem [285] : 
                        (N11)? \nz.mem [382] : 1'b0;
  assign r_data_o[90] = (N8)? \nz.mem [90] : 
                        (N10)? \nz.mem [187] : 
                        (N9)? \nz.mem [284] : 
                        (N11)? \nz.mem [381] : 1'b0;
  assign r_data_o[89] = (N8)? \nz.mem [89] : 
                        (N10)? \nz.mem [186] : 
                        (N9)? \nz.mem [283] : 
                        (N11)? \nz.mem [380] : 1'b0;
  assign r_data_o[88] = (N8)? \nz.mem [88] : 
                        (N10)? \nz.mem [185] : 
                        (N9)? \nz.mem [282] : 
                        (N11)? \nz.mem [379] : 1'b0;
  assign r_data_o[87] = (N8)? \nz.mem [87] : 
                        (N10)? \nz.mem [184] : 
                        (N9)? \nz.mem [281] : 
                        (N11)? \nz.mem [378] : 1'b0;
  assign r_data_o[86] = (N8)? \nz.mem [86] : 
                        (N10)? \nz.mem [183] : 
                        (N9)? \nz.mem [280] : 
                        (N11)? \nz.mem [377] : 1'b0;
  assign r_data_o[85] = (N8)? \nz.mem [85] : 
                        (N10)? \nz.mem [182] : 
                        (N9)? \nz.mem [279] : 
                        (N11)? \nz.mem [376] : 1'b0;
  assign r_data_o[84] = (N8)? \nz.mem [84] : 
                        (N10)? \nz.mem [181] : 
                        (N9)? \nz.mem [278] : 
                        (N11)? \nz.mem [375] : 1'b0;
  assign r_data_o[83] = (N8)? \nz.mem [83] : 
                        (N10)? \nz.mem [180] : 
                        (N9)? \nz.mem [277] : 
                        (N11)? \nz.mem [374] : 1'b0;
  assign r_data_o[82] = (N8)? \nz.mem [82] : 
                        (N10)? \nz.mem [179] : 
                        (N9)? \nz.mem [276] : 
                        (N11)? \nz.mem [373] : 1'b0;
  assign r_data_o[81] = (N8)? \nz.mem [81] : 
                        (N10)? \nz.mem [178] : 
                        (N9)? \nz.mem [275] : 
                        (N11)? \nz.mem [372] : 1'b0;
  assign r_data_o[80] = (N8)? \nz.mem [80] : 
                        (N10)? \nz.mem [177] : 
                        (N9)? \nz.mem [274] : 
                        (N11)? \nz.mem [371] : 1'b0;
  assign r_data_o[79] = (N8)? \nz.mem [79] : 
                        (N10)? \nz.mem [176] : 
                        (N9)? \nz.mem [273] : 
                        (N11)? \nz.mem [370] : 1'b0;
  assign r_data_o[78] = (N8)? \nz.mem [78] : 
                        (N10)? \nz.mem [175] : 
                        (N9)? \nz.mem [272] : 
                        (N11)? \nz.mem [369] : 1'b0;
  assign r_data_o[77] = (N8)? \nz.mem [77] : 
                        (N10)? \nz.mem [174] : 
                        (N9)? \nz.mem [271] : 
                        (N11)? \nz.mem [368] : 1'b0;
  assign r_data_o[76] = (N8)? \nz.mem [76] : 
                        (N10)? \nz.mem [173] : 
                        (N9)? \nz.mem [270] : 
                        (N11)? \nz.mem [367] : 1'b0;
  assign r_data_o[75] = (N8)? \nz.mem [75] : 
                        (N10)? \nz.mem [172] : 
                        (N9)? \nz.mem [269] : 
                        (N11)? \nz.mem [366] : 1'b0;
  assign r_data_o[74] = (N8)? \nz.mem [74] : 
                        (N10)? \nz.mem [171] : 
                        (N9)? \nz.mem [268] : 
                        (N11)? \nz.mem [365] : 1'b0;
  assign r_data_o[73] = (N8)? \nz.mem [73] : 
                        (N10)? \nz.mem [170] : 
                        (N9)? \nz.mem [267] : 
                        (N11)? \nz.mem [364] : 1'b0;
  assign r_data_o[72] = (N8)? \nz.mem [72] : 
                        (N10)? \nz.mem [169] : 
                        (N9)? \nz.mem [266] : 
                        (N11)? \nz.mem [363] : 1'b0;
  assign r_data_o[71] = (N8)? \nz.mem [71] : 
                        (N10)? \nz.mem [168] : 
                        (N9)? \nz.mem [265] : 
                        (N11)? \nz.mem [362] : 1'b0;
  assign r_data_o[70] = (N8)? \nz.mem [70] : 
                        (N10)? \nz.mem [167] : 
                        (N9)? \nz.mem [264] : 
                        (N11)? \nz.mem [361] : 1'b0;
  assign r_data_o[69] = (N8)? \nz.mem [69] : 
                        (N10)? \nz.mem [166] : 
                        (N9)? \nz.mem [263] : 
                        (N11)? \nz.mem [360] : 1'b0;
  assign r_data_o[68] = (N8)? \nz.mem [68] : 
                        (N10)? \nz.mem [165] : 
                        (N9)? \nz.mem [262] : 
                        (N11)? \nz.mem [359] : 1'b0;
  assign r_data_o[67] = (N8)? \nz.mem [67] : 
                        (N10)? \nz.mem [164] : 
                        (N9)? \nz.mem [261] : 
                        (N11)? \nz.mem [358] : 1'b0;
  assign r_data_o[66] = (N8)? \nz.mem [66] : 
                        (N10)? \nz.mem [163] : 
                        (N9)? \nz.mem [260] : 
                        (N11)? \nz.mem [357] : 1'b0;
  assign r_data_o[65] = (N8)? \nz.mem [65] : 
                        (N10)? \nz.mem [162] : 
                        (N9)? \nz.mem [259] : 
                        (N11)? \nz.mem [356] : 1'b0;
  assign r_data_o[64] = (N8)? \nz.mem [64] : 
                        (N10)? \nz.mem [161] : 
                        (N9)? \nz.mem [258] : 
                        (N11)? \nz.mem [355] : 1'b0;
  assign r_data_o[63] = (N8)? \nz.mem [63] : 
                        (N10)? \nz.mem [160] : 
                        (N9)? \nz.mem [257] : 
                        (N11)? \nz.mem [354] : 1'b0;
  assign r_data_o[62] = (N8)? \nz.mem [62] : 
                        (N10)? \nz.mem [159] : 
                        (N9)? \nz.mem [256] : 
                        (N11)? \nz.mem [353] : 1'b0;
  assign r_data_o[61] = (N8)? \nz.mem [61] : 
                        (N10)? \nz.mem [158] : 
                        (N9)? \nz.mem [255] : 
                        (N11)? \nz.mem [352] : 1'b0;
  assign r_data_o[60] = (N8)? \nz.mem [60] : 
                        (N10)? \nz.mem [157] : 
                        (N9)? \nz.mem [254] : 
                        (N11)? \nz.mem [351] : 1'b0;
  assign r_data_o[59] = (N8)? \nz.mem [59] : 
                        (N10)? \nz.mem [156] : 
                        (N9)? \nz.mem [253] : 
                        (N11)? \nz.mem [350] : 1'b0;
  assign r_data_o[58] = (N8)? \nz.mem [58] : 
                        (N10)? \nz.mem [155] : 
                        (N9)? \nz.mem [252] : 
                        (N11)? \nz.mem [349] : 1'b0;
  assign r_data_o[57] = (N8)? \nz.mem [57] : 
                        (N10)? \nz.mem [154] : 
                        (N9)? \nz.mem [251] : 
                        (N11)? \nz.mem [348] : 1'b0;
  assign r_data_o[56] = (N8)? \nz.mem [56] : 
                        (N10)? \nz.mem [153] : 
                        (N9)? \nz.mem [250] : 
                        (N11)? \nz.mem [347] : 1'b0;
  assign r_data_o[55] = (N8)? \nz.mem [55] : 
                        (N10)? \nz.mem [152] : 
                        (N9)? \nz.mem [249] : 
                        (N11)? \nz.mem [346] : 1'b0;
  assign r_data_o[54] = (N8)? \nz.mem [54] : 
                        (N10)? \nz.mem [151] : 
                        (N9)? \nz.mem [248] : 
                        (N11)? \nz.mem [345] : 1'b0;
  assign r_data_o[53] = (N8)? \nz.mem [53] : 
                        (N10)? \nz.mem [150] : 
                        (N9)? \nz.mem [247] : 
                        (N11)? \nz.mem [344] : 1'b0;
  assign r_data_o[52] = (N8)? \nz.mem [52] : 
                        (N10)? \nz.mem [149] : 
                        (N9)? \nz.mem [246] : 
                        (N11)? \nz.mem [343] : 1'b0;
  assign r_data_o[51] = (N8)? \nz.mem [51] : 
                        (N10)? \nz.mem [148] : 
                        (N9)? \nz.mem [245] : 
                        (N11)? \nz.mem [342] : 1'b0;
  assign r_data_o[50] = (N8)? \nz.mem [50] : 
                        (N10)? \nz.mem [147] : 
                        (N9)? \nz.mem [244] : 
                        (N11)? \nz.mem [341] : 1'b0;
  assign r_data_o[49] = (N8)? \nz.mem [49] : 
                        (N10)? \nz.mem [146] : 
                        (N9)? \nz.mem [243] : 
                        (N11)? \nz.mem [340] : 1'b0;
  assign r_data_o[48] = (N8)? \nz.mem [48] : 
                        (N10)? \nz.mem [145] : 
                        (N9)? \nz.mem [242] : 
                        (N11)? \nz.mem [339] : 1'b0;
  assign r_data_o[47] = (N8)? \nz.mem [47] : 
                        (N10)? \nz.mem [144] : 
                        (N9)? \nz.mem [241] : 
                        (N11)? \nz.mem [338] : 1'b0;
  assign r_data_o[46] = (N8)? \nz.mem [46] : 
                        (N10)? \nz.mem [143] : 
                        (N9)? \nz.mem [240] : 
                        (N11)? \nz.mem [337] : 1'b0;
  assign r_data_o[45] = (N8)? \nz.mem [45] : 
                        (N10)? \nz.mem [142] : 
                        (N9)? \nz.mem [239] : 
                        (N11)? \nz.mem [336] : 1'b0;
  assign r_data_o[44] = (N8)? \nz.mem [44] : 
                        (N10)? \nz.mem [141] : 
                        (N9)? \nz.mem [238] : 
                        (N11)? \nz.mem [335] : 1'b0;
  assign r_data_o[43] = (N8)? \nz.mem [43] : 
                        (N10)? \nz.mem [140] : 
                        (N9)? \nz.mem [237] : 
                        (N11)? \nz.mem [334] : 1'b0;
  assign r_data_o[42] = (N8)? \nz.mem [42] : 
                        (N10)? \nz.mem [139] : 
                        (N9)? \nz.mem [236] : 
                        (N11)? \nz.mem [333] : 1'b0;
  assign r_data_o[41] = (N8)? \nz.mem [41] : 
                        (N10)? \nz.mem [138] : 
                        (N9)? \nz.mem [235] : 
                        (N11)? \nz.mem [332] : 1'b0;
  assign r_data_o[40] = (N8)? \nz.mem [40] : 
                        (N10)? \nz.mem [137] : 
                        (N9)? \nz.mem [234] : 
                        (N11)? \nz.mem [331] : 1'b0;
  assign r_data_o[39] = (N8)? \nz.mem [39] : 
                        (N10)? \nz.mem [136] : 
                        (N9)? \nz.mem [233] : 
                        (N11)? \nz.mem [330] : 1'b0;
  assign r_data_o[38] = (N8)? \nz.mem [38] : 
                        (N10)? \nz.mem [135] : 
                        (N9)? \nz.mem [232] : 
                        (N11)? \nz.mem [329] : 1'b0;
  assign r_data_o[37] = (N8)? \nz.mem [37] : 
                        (N10)? \nz.mem [134] : 
                        (N9)? \nz.mem [231] : 
                        (N11)? \nz.mem [328] : 1'b0;
  assign r_data_o[36] = (N8)? \nz.mem [36] : 
                        (N10)? \nz.mem [133] : 
                        (N9)? \nz.mem [230] : 
                        (N11)? \nz.mem [327] : 1'b0;
  assign r_data_o[35] = (N8)? \nz.mem [35] : 
                        (N10)? \nz.mem [132] : 
                        (N9)? \nz.mem [229] : 
                        (N11)? \nz.mem [326] : 1'b0;
  assign r_data_o[34] = (N8)? \nz.mem [34] : 
                        (N10)? \nz.mem [131] : 
                        (N9)? \nz.mem [228] : 
                        (N11)? \nz.mem [325] : 1'b0;
  assign r_data_o[33] = (N8)? \nz.mem [33] : 
                        (N10)? \nz.mem [130] : 
                        (N9)? \nz.mem [227] : 
                        (N11)? \nz.mem [324] : 1'b0;
  assign r_data_o[32] = (N8)? \nz.mem [32] : 
                        (N10)? \nz.mem [129] : 
                        (N9)? \nz.mem [226] : 
                        (N11)? \nz.mem [323] : 1'b0;
  assign r_data_o[31] = (N8)? \nz.mem [31] : 
                        (N10)? \nz.mem [128] : 
                        (N9)? \nz.mem [225] : 
                        (N11)? \nz.mem [322] : 1'b0;
  assign r_data_o[30] = (N8)? \nz.mem [30] : 
                        (N10)? \nz.mem [127] : 
                        (N9)? \nz.mem [224] : 
                        (N11)? \nz.mem [321] : 1'b0;
  assign r_data_o[29] = (N8)? \nz.mem [29] : 
                        (N10)? \nz.mem [126] : 
                        (N9)? \nz.mem [223] : 
                        (N11)? \nz.mem [320] : 1'b0;
  assign r_data_o[28] = (N8)? \nz.mem [28] : 
                        (N10)? \nz.mem [125] : 
                        (N9)? \nz.mem [222] : 
                        (N11)? \nz.mem [319] : 1'b0;
  assign r_data_o[27] = (N8)? \nz.mem [27] : 
                        (N10)? \nz.mem [124] : 
                        (N9)? \nz.mem [221] : 
                        (N11)? \nz.mem [318] : 1'b0;
  assign r_data_o[26] = (N8)? \nz.mem [26] : 
                        (N10)? \nz.mem [123] : 
                        (N9)? \nz.mem [220] : 
                        (N11)? \nz.mem [317] : 1'b0;
  assign r_data_o[25] = (N8)? \nz.mem [25] : 
                        (N10)? \nz.mem [122] : 
                        (N9)? \nz.mem [219] : 
                        (N11)? \nz.mem [316] : 1'b0;
  assign r_data_o[24] = (N8)? \nz.mem [24] : 
                        (N10)? \nz.mem [121] : 
                        (N9)? \nz.mem [218] : 
                        (N11)? \nz.mem [315] : 1'b0;
  assign r_data_o[23] = (N8)? \nz.mem [23] : 
                        (N10)? \nz.mem [120] : 
                        (N9)? \nz.mem [217] : 
                        (N11)? \nz.mem [314] : 1'b0;
  assign r_data_o[22] = (N8)? \nz.mem [22] : 
                        (N10)? \nz.mem [119] : 
                        (N9)? \nz.mem [216] : 
                        (N11)? \nz.mem [313] : 1'b0;
  assign r_data_o[21] = (N8)? \nz.mem [21] : 
                        (N10)? \nz.mem [118] : 
                        (N9)? \nz.mem [215] : 
                        (N11)? \nz.mem [312] : 1'b0;
  assign r_data_o[20] = (N8)? \nz.mem [20] : 
                        (N10)? \nz.mem [117] : 
                        (N9)? \nz.mem [214] : 
                        (N11)? \nz.mem [311] : 1'b0;
  assign r_data_o[19] = (N8)? \nz.mem [19] : 
                        (N10)? \nz.mem [116] : 
                        (N9)? \nz.mem [213] : 
                        (N11)? \nz.mem [310] : 1'b0;
  assign r_data_o[18] = (N8)? \nz.mem [18] : 
                        (N10)? \nz.mem [115] : 
                        (N9)? \nz.mem [212] : 
                        (N11)? \nz.mem [309] : 1'b0;
  assign r_data_o[17] = (N8)? \nz.mem [17] : 
                        (N10)? \nz.mem [114] : 
                        (N9)? \nz.mem [211] : 
                        (N11)? \nz.mem [308] : 1'b0;
  assign r_data_o[16] = (N8)? \nz.mem [16] : 
                        (N10)? \nz.mem [113] : 
                        (N9)? \nz.mem [210] : 
                        (N11)? \nz.mem [307] : 1'b0;
  assign r_data_o[15] = (N8)? \nz.mem [15] : 
                        (N10)? \nz.mem [112] : 
                        (N9)? \nz.mem [209] : 
                        (N11)? \nz.mem [306] : 1'b0;
  assign r_data_o[14] = (N8)? \nz.mem [14] : 
                        (N10)? \nz.mem [111] : 
                        (N9)? \nz.mem [208] : 
                        (N11)? \nz.mem [305] : 1'b0;
  assign r_data_o[13] = (N8)? \nz.mem [13] : 
                        (N10)? \nz.mem [110] : 
                        (N9)? \nz.mem [207] : 
                        (N11)? \nz.mem [304] : 1'b0;
  assign r_data_o[12] = (N8)? \nz.mem [12] : 
                        (N10)? \nz.mem [109] : 
                        (N9)? \nz.mem [206] : 
                        (N11)? \nz.mem [303] : 1'b0;
  assign r_data_o[11] = (N8)? \nz.mem [11] : 
                        (N10)? \nz.mem [108] : 
                        (N9)? \nz.mem [205] : 
                        (N11)? \nz.mem [302] : 1'b0;
  assign r_data_o[10] = (N8)? \nz.mem [10] : 
                        (N10)? \nz.mem [107] : 
                        (N9)? \nz.mem [204] : 
                        (N11)? \nz.mem [301] : 1'b0;
  assign r_data_o[9] = (N8)? \nz.mem [9] : 
                       (N10)? \nz.mem [106] : 
                       (N9)? \nz.mem [203] : 
                       (N11)? \nz.mem [300] : 1'b0;
  assign r_data_o[8] = (N8)? \nz.mem [8] : 
                       (N10)? \nz.mem [105] : 
                       (N9)? \nz.mem [202] : 
                       (N11)? \nz.mem [299] : 1'b0;
  assign r_data_o[7] = (N8)? \nz.mem [7] : 
                       (N10)? \nz.mem [104] : 
                       (N9)? \nz.mem [201] : 
                       (N11)? \nz.mem [298] : 1'b0;
  assign r_data_o[6] = (N8)? \nz.mem [6] : 
                       (N10)? \nz.mem [103] : 
                       (N9)? \nz.mem [200] : 
                       (N11)? \nz.mem [297] : 1'b0;
  assign r_data_o[5] = (N8)? \nz.mem [5] : 
                       (N10)? \nz.mem [102] : 
                       (N9)? \nz.mem [199] : 
                       (N11)? \nz.mem [296] : 1'b0;
  assign r_data_o[4] = (N8)? \nz.mem [4] : 
                       (N10)? \nz.mem [101] : 
                       (N9)? \nz.mem [198] : 
                       (N11)? \nz.mem [295] : 1'b0;
  assign r_data_o[3] = (N8)? \nz.mem [3] : 
                       (N10)? \nz.mem [100] : 
                       (N9)? \nz.mem [197] : 
                       (N11)? \nz.mem [294] : 1'b0;
  assign r_data_o[2] = (N8)? \nz.mem [2] : 
                       (N10)? \nz.mem [99] : 
                       (N9)? \nz.mem [196] : 
                       (N11)? \nz.mem [293] : 1'b0;
  assign r_data_o[1] = (N8)? \nz.mem [1] : 
                       (N10)? \nz.mem [98] : 
                       (N9)? \nz.mem [195] : 
                       (N11)? \nz.mem [292] : 1'b0;
  assign r_data_o[0] = (N8)? \nz.mem [0] : 
                       (N10)? \nz.mem [97] : 
                       (N9)? \nz.mem [194] : 
                       (N11)? \nz.mem [291] : 1'b0;
  assign N16 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign { N20, N19, N18, N17 } = (N4)? { N16, N15, N14, N13 } : 
                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = w_v_i;
  assign N5 = N12;
  assign N6 = ~r_addr_i[0];
  assign N7 = ~r_addr_i[1];
  assign N8 = N6 & N7;
  assign N9 = N6 & r_addr_i[1];
  assign N10 = r_addr_i[0] & N7;
  assign N11 = r_addr_i[0] & r_addr_i[1];
  assign N12 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N20) begin
      \nz.mem_387_sv2v_reg  <= w_data_i[96];
      \nz.mem_386_sv2v_reg  <= w_data_i[95];
      \nz.mem_385_sv2v_reg  <= w_data_i[94];
      \nz.mem_384_sv2v_reg  <= w_data_i[93];
      \nz.mem_383_sv2v_reg  <= w_data_i[92];
      \nz.mem_382_sv2v_reg  <= w_data_i[91];
      \nz.mem_381_sv2v_reg  <= w_data_i[90];
      \nz.mem_380_sv2v_reg  <= w_data_i[89];
      \nz.mem_379_sv2v_reg  <= w_data_i[88];
      \nz.mem_378_sv2v_reg  <= w_data_i[87];
      \nz.mem_377_sv2v_reg  <= w_data_i[86];
      \nz.mem_376_sv2v_reg  <= w_data_i[85];
      \nz.mem_375_sv2v_reg  <= w_data_i[84];
      \nz.mem_374_sv2v_reg  <= w_data_i[83];
      \nz.mem_373_sv2v_reg  <= w_data_i[82];
      \nz.mem_372_sv2v_reg  <= w_data_i[81];
      \nz.mem_371_sv2v_reg  <= w_data_i[80];
      \nz.mem_370_sv2v_reg  <= w_data_i[79];
      \nz.mem_369_sv2v_reg  <= w_data_i[78];
      \nz.mem_368_sv2v_reg  <= w_data_i[77];
      \nz.mem_367_sv2v_reg  <= w_data_i[76];
      \nz.mem_366_sv2v_reg  <= w_data_i[75];
      \nz.mem_365_sv2v_reg  <= w_data_i[74];
      \nz.mem_364_sv2v_reg  <= w_data_i[73];
      \nz.mem_363_sv2v_reg  <= w_data_i[72];
      \nz.mem_362_sv2v_reg  <= w_data_i[71];
      \nz.mem_361_sv2v_reg  <= w_data_i[70];
      \nz.mem_360_sv2v_reg  <= w_data_i[69];
      \nz.mem_359_sv2v_reg  <= w_data_i[68];
      \nz.mem_358_sv2v_reg  <= w_data_i[67];
      \nz.mem_357_sv2v_reg  <= w_data_i[66];
      \nz.mem_356_sv2v_reg  <= w_data_i[65];
      \nz.mem_355_sv2v_reg  <= w_data_i[64];
      \nz.mem_354_sv2v_reg  <= w_data_i[63];
      \nz.mem_353_sv2v_reg  <= w_data_i[62];
      \nz.mem_352_sv2v_reg  <= w_data_i[61];
      \nz.mem_351_sv2v_reg  <= w_data_i[60];
      \nz.mem_350_sv2v_reg  <= w_data_i[59];
      \nz.mem_349_sv2v_reg  <= w_data_i[58];
      \nz.mem_348_sv2v_reg  <= w_data_i[57];
      \nz.mem_347_sv2v_reg  <= w_data_i[56];
      \nz.mem_346_sv2v_reg  <= w_data_i[55];
      \nz.mem_345_sv2v_reg  <= w_data_i[54];
      \nz.mem_344_sv2v_reg  <= w_data_i[53];
      \nz.mem_343_sv2v_reg  <= w_data_i[52];
      \nz.mem_342_sv2v_reg  <= w_data_i[51];
      \nz.mem_341_sv2v_reg  <= w_data_i[50];
      \nz.mem_340_sv2v_reg  <= w_data_i[49];
      \nz.mem_339_sv2v_reg  <= w_data_i[48];
      \nz.mem_338_sv2v_reg  <= w_data_i[47];
      \nz.mem_337_sv2v_reg  <= w_data_i[46];
      \nz.mem_336_sv2v_reg  <= w_data_i[45];
      \nz.mem_335_sv2v_reg  <= w_data_i[44];
      \nz.mem_334_sv2v_reg  <= w_data_i[43];
      \nz.mem_333_sv2v_reg  <= w_data_i[42];
      \nz.mem_332_sv2v_reg  <= w_data_i[41];
      \nz.mem_331_sv2v_reg  <= w_data_i[40];
      \nz.mem_330_sv2v_reg  <= w_data_i[39];
      \nz.mem_329_sv2v_reg  <= w_data_i[38];
      \nz.mem_328_sv2v_reg  <= w_data_i[37];
      \nz.mem_327_sv2v_reg  <= w_data_i[36];
      \nz.mem_326_sv2v_reg  <= w_data_i[35];
      \nz.mem_325_sv2v_reg  <= w_data_i[34];
      \nz.mem_324_sv2v_reg  <= w_data_i[33];
      \nz.mem_323_sv2v_reg  <= w_data_i[32];
      \nz.mem_322_sv2v_reg  <= w_data_i[31];
      \nz.mem_321_sv2v_reg  <= w_data_i[30];
      \nz.mem_320_sv2v_reg  <= w_data_i[29];
      \nz.mem_319_sv2v_reg  <= w_data_i[28];
      \nz.mem_318_sv2v_reg  <= w_data_i[27];
      \nz.mem_317_sv2v_reg  <= w_data_i[26];
      \nz.mem_316_sv2v_reg  <= w_data_i[25];
      \nz.mem_315_sv2v_reg  <= w_data_i[24];
      \nz.mem_314_sv2v_reg  <= w_data_i[23];
      \nz.mem_313_sv2v_reg  <= w_data_i[22];
      \nz.mem_312_sv2v_reg  <= w_data_i[21];
      \nz.mem_311_sv2v_reg  <= w_data_i[20];
      \nz.mem_310_sv2v_reg  <= w_data_i[19];
      \nz.mem_309_sv2v_reg  <= w_data_i[18];
      \nz.mem_308_sv2v_reg  <= w_data_i[17];
      \nz.mem_307_sv2v_reg  <= w_data_i[16];
      \nz.mem_306_sv2v_reg  <= w_data_i[15];
      \nz.mem_305_sv2v_reg  <= w_data_i[14];
      \nz.mem_304_sv2v_reg  <= w_data_i[13];
      \nz.mem_303_sv2v_reg  <= w_data_i[12];
      \nz.mem_302_sv2v_reg  <= w_data_i[11];
      \nz.mem_301_sv2v_reg  <= w_data_i[10];
      \nz.mem_300_sv2v_reg  <= w_data_i[9];
      \nz.mem_299_sv2v_reg  <= w_data_i[8];
      \nz.mem_298_sv2v_reg  <= w_data_i[7];
      \nz.mem_297_sv2v_reg  <= w_data_i[6];
      \nz.mem_296_sv2v_reg  <= w_data_i[5];
      \nz.mem_295_sv2v_reg  <= w_data_i[4];
      \nz.mem_294_sv2v_reg  <= w_data_i[3];
      \nz.mem_293_sv2v_reg  <= w_data_i[2];
      \nz.mem_292_sv2v_reg  <= w_data_i[1];
      \nz.mem_291_sv2v_reg  <= w_data_i[0];
    end 
    if(N19) begin
      \nz.mem_290_sv2v_reg  <= w_data_i[96];
      \nz.mem_289_sv2v_reg  <= w_data_i[95];
      \nz.mem_288_sv2v_reg  <= w_data_i[94];
      \nz.mem_287_sv2v_reg  <= w_data_i[93];
      \nz.mem_286_sv2v_reg  <= w_data_i[92];
      \nz.mem_285_sv2v_reg  <= w_data_i[91];
      \nz.mem_284_sv2v_reg  <= w_data_i[90];
      \nz.mem_283_sv2v_reg  <= w_data_i[89];
      \nz.mem_282_sv2v_reg  <= w_data_i[88];
      \nz.mem_281_sv2v_reg  <= w_data_i[87];
      \nz.mem_280_sv2v_reg  <= w_data_i[86];
      \nz.mem_279_sv2v_reg  <= w_data_i[85];
      \nz.mem_278_sv2v_reg  <= w_data_i[84];
      \nz.mem_277_sv2v_reg  <= w_data_i[83];
      \nz.mem_276_sv2v_reg  <= w_data_i[82];
      \nz.mem_275_sv2v_reg  <= w_data_i[81];
      \nz.mem_274_sv2v_reg  <= w_data_i[80];
      \nz.mem_273_sv2v_reg  <= w_data_i[79];
      \nz.mem_272_sv2v_reg  <= w_data_i[78];
      \nz.mem_271_sv2v_reg  <= w_data_i[77];
      \nz.mem_270_sv2v_reg  <= w_data_i[76];
      \nz.mem_269_sv2v_reg  <= w_data_i[75];
      \nz.mem_268_sv2v_reg  <= w_data_i[74];
      \nz.mem_267_sv2v_reg  <= w_data_i[73];
      \nz.mem_266_sv2v_reg  <= w_data_i[72];
      \nz.mem_265_sv2v_reg  <= w_data_i[71];
      \nz.mem_264_sv2v_reg  <= w_data_i[70];
      \nz.mem_263_sv2v_reg  <= w_data_i[69];
      \nz.mem_262_sv2v_reg  <= w_data_i[68];
      \nz.mem_261_sv2v_reg  <= w_data_i[67];
      \nz.mem_260_sv2v_reg  <= w_data_i[66];
      \nz.mem_259_sv2v_reg  <= w_data_i[65];
      \nz.mem_258_sv2v_reg  <= w_data_i[64];
      \nz.mem_257_sv2v_reg  <= w_data_i[63];
      \nz.mem_256_sv2v_reg  <= w_data_i[62];
      \nz.mem_255_sv2v_reg  <= w_data_i[61];
      \nz.mem_254_sv2v_reg  <= w_data_i[60];
      \nz.mem_253_sv2v_reg  <= w_data_i[59];
      \nz.mem_252_sv2v_reg  <= w_data_i[58];
      \nz.mem_251_sv2v_reg  <= w_data_i[57];
      \nz.mem_250_sv2v_reg  <= w_data_i[56];
      \nz.mem_249_sv2v_reg  <= w_data_i[55];
      \nz.mem_248_sv2v_reg  <= w_data_i[54];
      \nz.mem_247_sv2v_reg  <= w_data_i[53];
      \nz.mem_246_sv2v_reg  <= w_data_i[52];
      \nz.mem_245_sv2v_reg  <= w_data_i[51];
      \nz.mem_244_sv2v_reg  <= w_data_i[50];
      \nz.mem_243_sv2v_reg  <= w_data_i[49];
      \nz.mem_242_sv2v_reg  <= w_data_i[48];
      \nz.mem_241_sv2v_reg  <= w_data_i[47];
      \nz.mem_240_sv2v_reg  <= w_data_i[46];
      \nz.mem_239_sv2v_reg  <= w_data_i[45];
      \nz.mem_238_sv2v_reg  <= w_data_i[44];
      \nz.mem_237_sv2v_reg  <= w_data_i[43];
      \nz.mem_236_sv2v_reg  <= w_data_i[42];
      \nz.mem_235_sv2v_reg  <= w_data_i[41];
      \nz.mem_234_sv2v_reg  <= w_data_i[40];
      \nz.mem_233_sv2v_reg  <= w_data_i[39];
      \nz.mem_232_sv2v_reg  <= w_data_i[38];
      \nz.mem_231_sv2v_reg  <= w_data_i[37];
      \nz.mem_230_sv2v_reg  <= w_data_i[36];
      \nz.mem_229_sv2v_reg  <= w_data_i[35];
      \nz.mem_228_sv2v_reg  <= w_data_i[34];
      \nz.mem_227_sv2v_reg  <= w_data_i[33];
      \nz.mem_226_sv2v_reg  <= w_data_i[32];
      \nz.mem_225_sv2v_reg  <= w_data_i[31];
      \nz.mem_224_sv2v_reg  <= w_data_i[30];
      \nz.mem_223_sv2v_reg  <= w_data_i[29];
      \nz.mem_222_sv2v_reg  <= w_data_i[28];
      \nz.mem_221_sv2v_reg  <= w_data_i[27];
      \nz.mem_220_sv2v_reg  <= w_data_i[26];
      \nz.mem_219_sv2v_reg  <= w_data_i[25];
      \nz.mem_218_sv2v_reg  <= w_data_i[24];
      \nz.mem_217_sv2v_reg  <= w_data_i[23];
      \nz.mem_216_sv2v_reg  <= w_data_i[22];
      \nz.mem_215_sv2v_reg  <= w_data_i[21];
      \nz.mem_214_sv2v_reg  <= w_data_i[20];
      \nz.mem_213_sv2v_reg  <= w_data_i[19];
      \nz.mem_212_sv2v_reg  <= w_data_i[18];
      \nz.mem_211_sv2v_reg  <= w_data_i[17];
      \nz.mem_210_sv2v_reg  <= w_data_i[16];
      \nz.mem_209_sv2v_reg  <= w_data_i[15];
      \nz.mem_208_sv2v_reg  <= w_data_i[14];
      \nz.mem_207_sv2v_reg  <= w_data_i[13];
      \nz.mem_206_sv2v_reg  <= w_data_i[12];
      \nz.mem_205_sv2v_reg  <= w_data_i[11];
      \nz.mem_204_sv2v_reg  <= w_data_i[10];
      \nz.mem_203_sv2v_reg  <= w_data_i[9];
      \nz.mem_202_sv2v_reg  <= w_data_i[8];
      \nz.mem_201_sv2v_reg  <= w_data_i[7];
      \nz.mem_200_sv2v_reg  <= w_data_i[6];
      \nz.mem_199_sv2v_reg  <= w_data_i[5];
      \nz.mem_198_sv2v_reg  <= w_data_i[4];
      \nz.mem_197_sv2v_reg  <= w_data_i[3];
      \nz.mem_196_sv2v_reg  <= w_data_i[2];
      \nz.mem_195_sv2v_reg  <= w_data_i[1];
      \nz.mem_194_sv2v_reg  <= w_data_i[0];
    end 
    if(N18) begin
      \nz.mem_193_sv2v_reg  <= w_data_i[96];
      \nz.mem_192_sv2v_reg  <= w_data_i[95];
      \nz.mem_191_sv2v_reg  <= w_data_i[94];
      \nz.mem_190_sv2v_reg  <= w_data_i[93];
      \nz.mem_189_sv2v_reg  <= w_data_i[92];
      \nz.mem_188_sv2v_reg  <= w_data_i[91];
      \nz.mem_187_sv2v_reg  <= w_data_i[90];
      \nz.mem_186_sv2v_reg  <= w_data_i[89];
      \nz.mem_185_sv2v_reg  <= w_data_i[88];
      \nz.mem_184_sv2v_reg  <= w_data_i[87];
      \nz.mem_183_sv2v_reg  <= w_data_i[86];
      \nz.mem_182_sv2v_reg  <= w_data_i[85];
      \nz.mem_181_sv2v_reg  <= w_data_i[84];
      \nz.mem_180_sv2v_reg  <= w_data_i[83];
      \nz.mem_179_sv2v_reg  <= w_data_i[82];
      \nz.mem_178_sv2v_reg  <= w_data_i[81];
      \nz.mem_177_sv2v_reg  <= w_data_i[80];
      \nz.mem_176_sv2v_reg  <= w_data_i[79];
      \nz.mem_175_sv2v_reg  <= w_data_i[78];
      \nz.mem_174_sv2v_reg  <= w_data_i[77];
      \nz.mem_173_sv2v_reg  <= w_data_i[76];
      \nz.mem_172_sv2v_reg  <= w_data_i[75];
      \nz.mem_171_sv2v_reg  <= w_data_i[74];
      \nz.mem_170_sv2v_reg  <= w_data_i[73];
      \nz.mem_169_sv2v_reg  <= w_data_i[72];
      \nz.mem_168_sv2v_reg  <= w_data_i[71];
      \nz.mem_167_sv2v_reg  <= w_data_i[70];
      \nz.mem_166_sv2v_reg  <= w_data_i[69];
      \nz.mem_165_sv2v_reg  <= w_data_i[68];
      \nz.mem_164_sv2v_reg  <= w_data_i[67];
      \nz.mem_163_sv2v_reg  <= w_data_i[66];
      \nz.mem_162_sv2v_reg  <= w_data_i[65];
      \nz.mem_161_sv2v_reg  <= w_data_i[64];
      \nz.mem_160_sv2v_reg  <= w_data_i[63];
      \nz.mem_159_sv2v_reg  <= w_data_i[62];
      \nz.mem_158_sv2v_reg  <= w_data_i[61];
      \nz.mem_157_sv2v_reg  <= w_data_i[60];
      \nz.mem_156_sv2v_reg  <= w_data_i[59];
      \nz.mem_155_sv2v_reg  <= w_data_i[58];
      \nz.mem_154_sv2v_reg  <= w_data_i[57];
      \nz.mem_153_sv2v_reg  <= w_data_i[56];
      \nz.mem_152_sv2v_reg  <= w_data_i[55];
      \nz.mem_151_sv2v_reg  <= w_data_i[54];
      \nz.mem_150_sv2v_reg  <= w_data_i[53];
      \nz.mem_149_sv2v_reg  <= w_data_i[52];
      \nz.mem_148_sv2v_reg  <= w_data_i[51];
      \nz.mem_147_sv2v_reg  <= w_data_i[50];
      \nz.mem_146_sv2v_reg  <= w_data_i[49];
      \nz.mem_145_sv2v_reg  <= w_data_i[48];
      \nz.mem_144_sv2v_reg  <= w_data_i[47];
      \nz.mem_143_sv2v_reg  <= w_data_i[46];
      \nz.mem_142_sv2v_reg  <= w_data_i[45];
      \nz.mem_141_sv2v_reg  <= w_data_i[44];
      \nz.mem_140_sv2v_reg  <= w_data_i[43];
      \nz.mem_139_sv2v_reg  <= w_data_i[42];
      \nz.mem_138_sv2v_reg  <= w_data_i[41];
      \nz.mem_137_sv2v_reg  <= w_data_i[40];
      \nz.mem_136_sv2v_reg  <= w_data_i[39];
      \nz.mem_135_sv2v_reg  <= w_data_i[38];
      \nz.mem_134_sv2v_reg  <= w_data_i[37];
      \nz.mem_133_sv2v_reg  <= w_data_i[36];
      \nz.mem_132_sv2v_reg  <= w_data_i[35];
      \nz.mem_131_sv2v_reg  <= w_data_i[34];
      \nz.mem_130_sv2v_reg  <= w_data_i[33];
      \nz.mem_129_sv2v_reg  <= w_data_i[32];
      \nz.mem_128_sv2v_reg  <= w_data_i[31];
      \nz.mem_127_sv2v_reg  <= w_data_i[30];
      \nz.mem_126_sv2v_reg  <= w_data_i[29];
      \nz.mem_125_sv2v_reg  <= w_data_i[28];
      \nz.mem_124_sv2v_reg  <= w_data_i[27];
      \nz.mem_123_sv2v_reg  <= w_data_i[26];
      \nz.mem_122_sv2v_reg  <= w_data_i[25];
      \nz.mem_121_sv2v_reg  <= w_data_i[24];
      \nz.mem_120_sv2v_reg  <= w_data_i[23];
      \nz.mem_119_sv2v_reg  <= w_data_i[22];
      \nz.mem_118_sv2v_reg  <= w_data_i[21];
      \nz.mem_117_sv2v_reg  <= w_data_i[20];
      \nz.mem_116_sv2v_reg  <= w_data_i[19];
      \nz.mem_115_sv2v_reg  <= w_data_i[18];
      \nz.mem_114_sv2v_reg  <= w_data_i[17];
      \nz.mem_113_sv2v_reg  <= w_data_i[16];
      \nz.mem_112_sv2v_reg  <= w_data_i[15];
      \nz.mem_111_sv2v_reg  <= w_data_i[14];
      \nz.mem_110_sv2v_reg  <= w_data_i[13];
      \nz.mem_109_sv2v_reg  <= w_data_i[12];
      \nz.mem_108_sv2v_reg  <= w_data_i[11];
      \nz.mem_107_sv2v_reg  <= w_data_i[10];
      \nz.mem_106_sv2v_reg  <= w_data_i[9];
      \nz.mem_105_sv2v_reg  <= w_data_i[8];
      \nz.mem_104_sv2v_reg  <= w_data_i[7];
      \nz.mem_103_sv2v_reg  <= w_data_i[6];
      \nz.mem_102_sv2v_reg  <= w_data_i[5];
      \nz.mem_101_sv2v_reg  <= w_data_i[4];
      \nz.mem_100_sv2v_reg  <= w_data_i[3];
      \nz.mem_99_sv2v_reg  <= w_data_i[2];
      \nz.mem_98_sv2v_reg  <= w_data_i[1];
      \nz.mem_97_sv2v_reg  <= w_data_i[0];
    end 
    if(N17) begin
      \nz.mem_96_sv2v_reg  <= w_data_i[96];
      \nz.mem_95_sv2v_reg  <= w_data_i[95];
      \nz.mem_94_sv2v_reg  <= w_data_i[94];
      \nz.mem_93_sv2v_reg  <= w_data_i[93];
      \nz.mem_92_sv2v_reg  <= w_data_i[92];
      \nz.mem_91_sv2v_reg  <= w_data_i[91];
      \nz.mem_90_sv2v_reg  <= w_data_i[90];
      \nz.mem_89_sv2v_reg  <= w_data_i[89];
      \nz.mem_88_sv2v_reg  <= w_data_i[88];
      \nz.mem_87_sv2v_reg  <= w_data_i[87];
      \nz.mem_86_sv2v_reg  <= w_data_i[86];
      \nz.mem_85_sv2v_reg  <= w_data_i[85];
      \nz.mem_84_sv2v_reg  <= w_data_i[84];
      \nz.mem_83_sv2v_reg  <= w_data_i[83];
      \nz.mem_82_sv2v_reg  <= w_data_i[82];
      \nz.mem_81_sv2v_reg  <= w_data_i[81];
      \nz.mem_80_sv2v_reg  <= w_data_i[80];
      \nz.mem_79_sv2v_reg  <= w_data_i[79];
      \nz.mem_78_sv2v_reg  <= w_data_i[78];
      \nz.mem_77_sv2v_reg  <= w_data_i[77];
      \nz.mem_76_sv2v_reg  <= w_data_i[76];
      \nz.mem_75_sv2v_reg  <= w_data_i[75];
      \nz.mem_74_sv2v_reg  <= w_data_i[74];
      \nz.mem_73_sv2v_reg  <= w_data_i[73];
      \nz.mem_72_sv2v_reg  <= w_data_i[72];
      \nz.mem_71_sv2v_reg  <= w_data_i[71];
      \nz.mem_70_sv2v_reg  <= w_data_i[70];
      \nz.mem_69_sv2v_reg  <= w_data_i[69];
      \nz.mem_68_sv2v_reg  <= w_data_i[68];
      \nz.mem_67_sv2v_reg  <= w_data_i[67];
      \nz.mem_66_sv2v_reg  <= w_data_i[66];
      \nz.mem_65_sv2v_reg  <= w_data_i[65];
      \nz.mem_64_sv2v_reg  <= w_data_i[64];
      \nz.mem_63_sv2v_reg  <= w_data_i[63];
      \nz.mem_62_sv2v_reg  <= w_data_i[62];
      \nz.mem_61_sv2v_reg  <= w_data_i[61];
      \nz.mem_60_sv2v_reg  <= w_data_i[60];
      \nz.mem_59_sv2v_reg  <= w_data_i[59];
      \nz.mem_58_sv2v_reg  <= w_data_i[58];
      \nz.mem_57_sv2v_reg  <= w_data_i[57];
      \nz.mem_56_sv2v_reg  <= w_data_i[56];
      \nz.mem_55_sv2v_reg  <= w_data_i[55];
      \nz.mem_54_sv2v_reg  <= w_data_i[54];
      \nz.mem_53_sv2v_reg  <= w_data_i[53];
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p97_els_p4_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [96:0] w_data_i;
  input [1:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;

  bsg_mem_1r1w_synth_width_p97_els_p4_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p97_els_p4_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [96:0] data_i;
  output [96:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [96:0] data_o;
  wire ready_o,v_o,enque,full,empty,sv2v_dc_1,sv2v_dc_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p4
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p97_els_p4_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_o;
  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p97_els_p4
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [96:0] data_i;
  output [96:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [96:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p97_els_p4_ready_THEN_valid_p0
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_mem_1r1w_synth_width_p53_els_p2_read_write_same_addr_p1_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [52:0] w_data_i;
  input [0:0] r_addr_i;
  output [52:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [52:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [105:0] \nz.mem ;
  reg \nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,
  \nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,
  \nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,
  \nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,
  \nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,
  \nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,
  \nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[52] = (N3)? \nz.mem [52] : 
                        (N0)? \nz.mem [105] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[51] = (N3)? \nz.mem [51] : 
                        (N0)? \nz.mem [104] : 1'b0;
  assign r_data_o[50] = (N3)? \nz.mem [50] : 
                        (N0)? \nz.mem [103] : 1'b0;
  assign r_data_o[49] = (N3)? \nz.mem [49] : 
                        (N0)? \nz.mem [102] : 1'b0;
  assign r_data_o[48] = (N3)? \nz.mem [48] : 
                        (N0)? \nz.mem [101] : 1'b0;
  assign r_data_o[47] = (N3)? \nz.mem [47] : 
                        (N0)? \nz.mem [100] : 1'b0;
  assign r_data_o[46] = (N3)? \nz.mem [46] : 
                        (N0)? \nz.mem [99] : 1'b0;
  assign r_data_o[45] = (N3)? \nz.mem [45] : 
                        (N0)? \nz.mem [98] : 1'b0;
  assign r_data_o[44] = (N3)? \nz.mem [44] : 
                        (N0)? \nz.mem [97] : 1'b0;
  assign r_data_o[43] = (N3)? \nz.mem [43] : 
                        (N0)? \nz.mem [96] : 1'b0;
  assign r_data_o[42] = (N3)? \nz.mem [42] : 
                        (N0)? \nz.mem [95] : 1'b0;
  assign r_data_o[41] = (N3)? \nz.mem [41] : 
                        (N0)? \nz.mem [94] : 1'b0;
  assign r_data_o[40] = (N3)? \nz.mem [40] : 
                        (N0)? \nz.mem [93] : 1'b0;
  assign r_data_o[39] = (N3)? \nz.mem [39] : 
                        (N0)? \nz.mem [92] : 1'b0;
  assign r_data_o[38] = (N3)? \nz.mem [38] : 
                        (N0)? \nz.mem [91] : 1'b0;
  assign r_data_o[37] = (N3)? \nz.mem [37] : 
                        (N0)? \nz.mem [90] : 1'b0;
  assign r_data_o[36] = (N3)? \nz.mem [36] : 
                        (N0)? \nz.mem [89] : 1'b0;
  assign r_data_o[35] = (N3)? \nz.mem [35] : 
                        (N0)? \nz.mem [88] : 1'b0;
  assign r_data_o[34] = (N3)? \nz.mem [34] : 
                        (N0)? \nz.mem [87] : 1'b0;
  assign r_data_o[33] = (N3)? \nz.mem [33] : 
                        (N0)? \nz.mem [86] : 1'b0;
  assign r_data_o[32] = (N3)? \nz.mem [32] : 
                        (N0)? \nz.mem [85] : 1'b0;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [84] : 1'b0;
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [83] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [82] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [81] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [80] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [79] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [78] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [77] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [76] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [75] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [74] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [73] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [72] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [71] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [70] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [69] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [68] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [67] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [66] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [65] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [64] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [63] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [62] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [61] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [60] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [59] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [58] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [57] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [56] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [55] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [54] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [53] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_105_sv2v_reg  <= w_data_i[52];
      \nz.mem_104_sv2v_reg  <= w_data_i[51];
      \nz.mem_103_sv2v_reg  <= w_data_i[50];
      \nz.mem_102_sv2v_reg  <= w_data_i[49];
      \nz.mem_101_sv2v_reg  <= w_data_i[48];
      \nz.mem_100_sv2v_reg  <= w_data_i[47];
      \nz.mem_99_sv2v_reg  <= w_data_i[46];
      \nz.mem_98_sv2v_reg  <= w_data_i[45];
      \nz.mem_97_sv2v_reg  <= w_data_i[44];
      \nz.mem_96_sv2v_reg  <= w_data_i[43];
      \nz.mem_95_sv2v_reg  <= w_data_i[42];
      \nz.mem_94_sv2v_reg  <= w_data_i[41];
      \nz.mem_93_sv2v_reg  <= w_data_i[40];
      \nz.mem_92_sv2v_reg  <= w_data_i[39];
      \nz.mem_91_sv2v_reg  <= w_data_i[38];
      \nz.mem_90_sv2v_reg  <= w_data_i[37];
      \nz.mem_89_sv2v_reg  <= w_data_i[36];
      \nz.mem_88_sv2v_reg  <= w_data_i[35];
      \nz.mem_87_sv2v_reg  <= w_data_i[34];
      \nz.mem_86_sv2v_reg  <= w_data_i[33];
      \nz.mem_85_sv2v_reg  <= w_data_i[32];
      \nz.mem_84_sv2v_reg  <= w_data_i[31];
      \nz.mem_83_sv2v_reg  <= w_data_i[30];
      \nz.mem_82_sv2v_reg  <= w_data_i[29];
      \nz.mem_81_sv2v_reg  <= w_data_i[28];
      \nz.mem_80_sv2v_reg  <= w_data_i[27];
      \nz.mem_79_sv2v_reg  <= w_data_i[26];
      \nz.mem_78_sv2v_reg  <= w_data_i[25];
      \nz.mem_77_sv2v_reg  <= w_data_i[24];
      \nz.mem_76_sv2v_reg  <= w_data_i[23];
      \nz.mem_75_sv2v_reg  <= w_data_i[22];
      \nz.mem_74_sv2v_reg  <= w_data_i[21];
      \nz.mem_73_sv2v_reg  <= w_data_i[20];
      \nz.mem_72_sv2v_reg  <= w_data_i[19];
      \nz.mem_71_sv2v_reg  <= w_data_i[18];
      \nz.mem_70_sv2v_reg  <= w_data_i[17];
      \nz.mem_69_sv2v_reg  <= w_data_i[16];
      \nz.mem_68_sv2v_reg  <= w_data_i[15];
      \nz.mem_67_sv2v_reg  <= w_data_i[14];
      \nz.mem_66_sv2v_reg  <= w_data_i[13];
      \nz.mem_65_sv2v_reg  <= w_data_i[12];
      \nz.mem_64_sv2v_reg  <= w_data_i[11];
      \nz.mem_63_sv2v_reg  <= w_data_i[10];
      \nz.mem_62_sv2v_reg  <= w_data_i[9];
      \nz.mem_61_sv2v_reg  <= w_data_i[8];
      \nz.mem_60_sv2v_reg  <= w_data_i[7];
      \nz.mem_59_sv2v_reg  <= w_data_i[6];
      \nz.mem_58_sv2v_reg  <= w_data_i[5];
      \nz.mem_57_sv2v_reg  <= w_data_i[4];
      \nz.mem_56_sv2v_reg  <= w_data_i[3];
      \nz.mem_55_sv2v_reg  <= w_data_i[2];
      \nz.mem_54_sv2v_reg  <= w_data_i[1];
      \nz.mem_53_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_52_sv2v_reg  <= w_data_i[52];
      \nz.mem_51_sv2v_reg  <= w_data_i[51];
      \nz.mem_50_sv2v_reg  <= w_data_i[50];
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p53_els_p2_read_write_same_addr_p1
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [52:0] w_data_i;
  input [0:0] r_addr_i;
  output [52:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [52:0] r_data_o;

  bsg_mem_1r1w_synth_width_p53_els_p2_read_write_same_addr_p1_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p53_allow_enq_deq_on_full_p1
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [52:0] data_i;
  output [52:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [52:0] data_o;
  wire ready_o,v_o,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,
  N10,N11,N12,N13,N14,N15,N16;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p53_els_p2_read_write_same_addr_p1
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign N1 = v_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N6 | N9;
  assign N6 = empty_r & N5;
  assign N5 = ~v_i;
  assign N9 = N8 & N5;
  assign N8 = N7 & yumi_i;
  assign N7 = ~full_r;
  assign N4 = N13 | N16;
  assign N13 = N11 & N12;
  assign N11 = N10 & v_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N16 = full_r & N15;
  assign N15 = ~N14;
  assign N14 = yumi_i ^ v_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_manycore_endpoint_x_cord_width_p7_y_cord_width_p7_fifo_els_p4_data_width_p32_addr_width_p28
(
  clk_i,
  reset_i,
  link_sif_i,
  link_sif_o,
  packet_o,
  packet_v_o,
  packet_yumi_i,
  return_packet_i,
  return_packet_v_i,
  return_packet_credit_or_ready_o,
  packet_i,
  packet_v_i,
  packet_credit_or_ready_o,
  return_packet_o,
  return_packet_v_o,
  return_packet_yumi_i,
  return_packet_fifo_full_o
);

  input [153:0] link_sif_i;
  output [153:0] link_sif_o;
  output [96:0] packet_o;
  input [52:0] return_packet_i;
  input [96:0] packet_i;
  output [52:0] return_packet_o;
  input clk_i;
  input reset_i;
  input packet_yumi_i;
  input return_packet_v_i;
  input packet_v_i;
  input return_packet_yumi_i;
  output packet_v_o;
  output return_packet_credit_or_ready_o;
  output packet_credit_or_ready_o;
  output return_packet_v_o;
  output return_packet_fifo_full_o;
  wire [153:0] link_sif_o;
  wire [96:0] packet_o;
  wire [52:0] return_packet_o;
  wire packet_v_o,return_packet_credit_or_ready_o,packet_credit_or_ready_o,
  return_packet_v_o,return_packet_fifo_full_o,link_sif_i_152_,link_sif_i_53_,link_sif_o_153_,
  link_sif_o_151_,link_sif_o_150_,link_sif_o_149_,link_sif_o_148_,link_sif_o_147_,
  link_sif_o_146_,link_sif_o_145_,link_sif_o_144_,link_sif_o_143_,link_sif_o_142_,
  link_sif_o_141_,link_sif_o_140_,link_sif_o_139_,link_sif_o_138_,link_sif_o_137_,
  link_sif_o_136_,link_sif_o_135_,link_sif_o_134_,link_sif_o_133_,link_sif_o_132_,
  link_sif_o_131_,link_sif_o_130_,link_sif_o_129_,link_sif_o_128_,link_sif_o_127_,
  link_sif_o_126_,link_sif_o_125_,link_sif_o_124_,link_sif_o_123_,link_sif_o_122_,
  link_sif_o_121_,link_sif_o_120_,link_sif_o_119_,link_sif_o_118_,link_sif_o_117_,
  link_sif_o_116_,link_sif_o_115_,link_sif_o_114_,link_sif_o_113_,link_sif_o_112_,
  link_sif_o_111_,link_sif_o_110_,link_sif_o_109_,link_sif_o_108_,link_sif_o_107_,
  link_sif_o_106_,link_sif_o_105_,link_sif_o_104_,link_sif_o_103_,link_sif_o_102_,
  link_sif_o_101_,link_sif_o_100_,link_sif_o_99_,link_sif_o_98_,link_sif_o_97_,
  link_sif_o_96_,link_sif_o_95_,link_sif_o_94_,link_sif_o_93_,link_sif_o_92_,
  link_sif_o_91_,link_sif_o_90_,link_sif_o_89_,link_sif_o_88_,link_sif_o_87_,
  link_sif_o_86_,link_sif_o_85_,link_sif_o_84_,link_sif_o_83_,link_sif_o_82_,link_sif_o_81_,
  link_sif_o_80_,link_sif_o_79_,link_sif_o_78_,link_sif_o_77_,link_sif_o_76_,
  link_sif_o_75_,link_sif_o_74_,link_sif_o_73_,link_sif_o_72_,link_sif_o_71_,
  link_sif_o_70_,link_sif_o_69_,link_sif_o_68_,link_sif_o_67_,link_sif_o_66_,link_sif_o_65_,
  link_sif_o_64_,link_sif_o_63_,link_sif_o_62_,link_sif_o_61_,link_sif_o_60_,
  link_sif_o_59_,link_sif_o_58_,link_sif_o_57_,link_sif_o_56_,link_sif_o_55_,
  link_sif_o_54_,link_sif_o_52_,link_sif_o_51_,link_sif_o_50_,link_sif_o_49_,link_sif_o_48_,
  link_sif_o_47_,link_sif_o_46_,link_sif_o_45_,link_sif_o_44_,link_sif_o_43_,
  link_sif_o_42_,link_sif_o_41_,link_sif_o_40_,link_sif_o_39_,link_sif_o_38_,
  link_sif_o_37_,link_sif_o_36_,link_sif_o_35_,link_sif_o_34_,link_sif_o_33_,link_sif_o_32_,
  link_sif_o_31_,link_sif_o_30_,link_sif_o_29_,link_sif_o_28_,link_sif_o_27_,
  link_sif_o_26_,link_sif_o_25_,link_sif_o_24_,link_sif_o_23_,link_sif_o_22_,
  link_sif_o_21_,link_sif_o_20_,link_sif_o_19_,link_sif_o_18_,link_sif_o_17_,link_sif_o_16_,
  link_sif_o_15_,link_sif_o_14_,link_sif_o_13_,link_sif_o_12_,link_sif_o_11_,
  link_sif_o_10_,link_sif_o_9_,link_sif_o_8_,link_sif_o_7_,link_sif_o_6_,link_sif_o_5_,
  link_sif_o_4_,link_sif_o_3_,link_sif_o_2_,link_sif_o_1_,link_sif_o_0_,
  returned_fifo_ready;
  assign link_sif_o[53] = 1'b1;
  assign link_sif_i_152_ = link_sif_i[152];
  assign packet_credit_or_ready_o = link_sif_i_152_;
  assign link_sif_i_53_ = link_sif_i[53];
  assign return_packet_credit_or_ready_o = link_sif_i_53_;
  assign link_sif_o_153_ = packet_v_i;
  assign link_sif_o[153] = link_sif_o_153_;
  assign link_sif_o_151_ = packet_i[96];
  assign link_sif_o[151] = link_sif_o_151_;
  assign link_sif_o_150_ = packet_i[95];
  assign link_sif_o[150] = link_sif_o_150_;
  assign link_sif_o_149_ = packet_i[94];
  assign link_sif_o[149] = link_sif_o_149_;
  assign link_sif_o_148_ = packet_i[93];
  assign link_sif_o[148] = link_sif_o_148_;
  assign link_sif_o_147_ = packet_i[92];
  assign link_sif_o[147] = link_sif_o_147_;
  assign link_sif_o_146_ = packet_i[91];
  assign link_sif_o[146] = link_sif_o_146_;
  assign link_sif_o_145_ = packet_i[90];
  assign link_sif_o[145] = link_sif_o_145_;
  assign link_sif_o_144_ = packet_i[89];
  assign link_sif_o[144] = link_sif_o_144_;
  assign link_sif_o_143_ = packet_i[88];
  assign link_sif_o[143] = link_sif_o_143_;
  assign link_sif_o_142_ = packet_i[87];
  assign link_sif_o[142] = link_sif_o_142_;
  assign link_sif_o_141_ = packet_i[86];
  assign link_sif_o[141] = link_sif_o_141_;
  assign link_sif_o_140_ = packet_i[85];
  assign link_sif_o[140] = link_sif_o_140_;
  assign link_sif_o_139_ = packet_i[84];
  assign link_sif_o[139] = link_sif_o_139_;
  assign link_sif_o_138_ = packet_i[83];
  assign link_sif_o[138] = link_sif_o_138_;
  assign link_sif_o_137_ = packet_i[82];
  assign link_sif_o[137] = link_sif_o_137_;
  assign link_sif_o_136_ = packet_i[81];
  assign link_sif_o[136] = link_sif_o_136_;
  assign link_sif_o_135_ = packet_i[80];
  assign link_sif_o[135] = link_sif_o_135_;
  assign link_sif_o_134_ = packet_i[79];
  assign link_sif_o[134] = link_sif_o_134_;
  assign link_sif_o_133_ = packet_i[78];
  assign link_sif_o[133] = link_sif_o_133_;
  assign link_sif_o_132_ = packet_i[77];
  assign link_sif_o[132] = link_sif_o_132_;
  assign link_sif_o_131_ = packet_i[76];
  assign link_sif_o[131] = link_sif_o_131_;
  assign link_sif_o_130_ = packet_i[75];
  assign link_sif_o[130] = link_sif_o_130_;
  assign link_sif_o_129_ = packet_i[74];
  assign link_sif_o[129] = link_sif_o_129_;
  assign link_sif_o_128_ = packet_i[73];
  assign link_sif_o[128] = link_sif_o_128_;
  assign link_sif_o_127_ = packet_i[72];
  assign link_sif_o[127] = link_sif_o_127_;
  assign link_sif_o_126_ = packet_i[71];
  assign link_sif_o[126] = link_sif_o_126_;
  assign link_sif_o_125_ = packet_i[70];
  assign link_sif_o[125] = link_sif_o_125_;
  assign link_sif_o_124_ = packet_i[69];
  assign link_sif_o[124] = link_sif_o_124_;
  assign link_sif_o_123_ = packet_i[68];
  assign link_sif_o[123] = link_sif_o_123_;
  assign link_sif_o_122_ = packet_i[67];
  assign link_sif_o[122] = link_sif_o_122_;
  assign link_sif_o_121_ = packet_i[66];
  assign link_sif_o[121] = link_sif_o_121_;
  assign link_sif_o_120_ = packet_i[65];
  assign link_sif_o[120] = link_sif_o_120_;
  assign link_sif_o_119_ = packet_i[64];
  assign link_sif_o[119] = link_sif_o_119_;
  assign link_sif_o_118_ = packet_i[63];
  assign link_sif_o[118] = link_sif_o_118_;
  assign link_sif_o_117_ = packet_i[62];
  assign link_sif_o[117] = link_sif_o_117_;
  assign link_sif_o_116_ = packet_i[61];
  assign link_sif_o[116] = link_sif_o_116_;
  assign link_sif_o_115_ = packet_i[60];
  assign link_sif_o[115] = link_sif_o_115_;
  assign link_sif_o_114_ = packet_i[59];
  assign link_sif_o[114] = link_sif_o_114_;
  assign link_sif_o_113_ = packet_i[58];
  assign link_sif_o[113] = link_sif_o_113_;
  assign link_sif_o_112_ = packet_i[57];
  assign link_sif_o[112] = link_sif_o_112_;
  assign link_sif_o_111_ = packet_i[56];
  assign link_sif_o[111] = link_sif_o_111_;
  assign link_sif_o_110_ = packet_i[55];
  assign link_sif_o[110] = link_sif_o_110_;
  assign link_sif_o_109_ = packet_i[54];
  assign link_sif_o[109] = link_sif_o_109_;
  assign link_sif_o_108_ = packet_i[53];
  assign link_sif_o[108] = link_sif_o_108_;
  assign link_sif_o_107_ = packet_i[52];
  assign link_sif_o[107] = link_sif_o_107_;
  assign link_sif_o_106_ = packet_i[51];
  assign link_sif_o[106] = link_sif_o_106_;
  assign link_sif_o_105_ = packet_i[50];
  assign link_sif_o[105] = link_sif_o_105_;
  assign link_sif_o_104_ = packet_i[49];
  assign link_sif_o[104] = link_sif_o_104_;
  assign link_sif_o_103_ = packet_i[48];
  assign link_sif_o[103] = link_sif_o_103_;
  assign link_sif_o_102_ = packet_i[47];
  assign link_sif_o[102] = link_sif_o_102_;
  assign link_sif_o_101_ = packet_i[46];
  assign link_sif_o[101] = link_sif_o_101_;
  assign link_sif_o_100_ = packet_i[45];
  assign link_sif_o[100] = link_sif_o_100_;
  assign link_sif_o_99_ = packet_i[44];
  assign link_sif_o[99] = link_sif_o_99_;
  assign link_sif_o_98_ = packet_i[43];
  assign link_sif_o[98] = link_sif_o_98_;
  assign link_sif_o_97_ = packet_i[42];
  assign link_sif_o[97] = link_sif_o_97_;
  assign link_sif_o_96_ = packet_i[41];
  assign link_sif_o[96] = link_sif_o_96_;
  assign link_sif_o_95_ = packet_i[40];
  assign link_sif_o[95] = link_sif_o_95_;
  assign link_sif_o_94_ = packet_i[39];
  assign link_sif_o[94] = link_sif_o_94_;
  assign link_sif_o_93_ = packet_i[38];
  assign link_sif_o[93] = link_sif_o_93_;
  assign link_sif_o_92_ = packet_i[37];
  assign link_sif_o[92] = link_sif_o_92_;
  assign link_sif_o_91_ = packet_i[36];
  assign link_sif_o[91] = link_sif_o_91_;
  assign link_sif_o_90_ = packet_i[35];
  assign link_sif_o[90] = link_sif_o_90_;
  assign link_sif_o_89_ = packet_i[34];
  assign link_sif_o[89] = link_sif_o_89_;
  assign link_sif_o_88_ = packet_i[33];
  assign link_sif_o[88] = link_sif_o_88_;
  assign link_sif_o_87_ = packet_i[32];
  assign link_sif_o[87] = link_sif_o_87_;
  assign link_sif_o_86_ = packet_i[31];
  assign link_sif_o[86] = link_sif_o_86_;
  assign link_sif_o_85_ = packet_i[30];
  assign link_sif_o[85] = link_sif_o_85_;
  assign link_sif_o_84_ = packet_i[29];
  assign link_sif_o[84] = link_sif_o_84_;
  assign link_sif_o_83_ = packet_i[28];
  assign link_sif_o[83] = link_sif_o_83_;
  assign link_sif_o_82_ = packet_i[27];
  assign link_sif_o[82] = link_sif_o_82_;
  assign link_sif_o_81_ = packet_i[26];
  assign link_sif_o[81] = link_sif_o_81_;
  assign link_sif_o_80_ = packet_i[25];
  assign link_sif_o[80] = link_sif_o_80_;
  assign link_sif_o_79_ = packet_i[24];
  assign link_sif_o[79] = link_sif_o_79_;
  assign link_sif_o_78_ = packet_i[23];
  assign link_sif_o[78] = link_sif_o_78_;
  assign link_sif_o_77_ = packet_i[22];
  assign link_sif_o[77] = link_sif_o_77_;
  assign link_sif_o_76_ = packet_i[21];
  assign link_sif_o[76] = link_sif_o_76_;
  assign link_sif_o_75_ = packet_i[20];
  assign link_sif_o[75] = link_sif_o_75_;
  assign link_sif_o_74_ = packet_i[19];
  assign link_sif_o[74] = link_sif_o_74_;
  assign link_sif_o_73_ = packet_i[18];
  assign link_sif_o[73] = link_sif_o_73_;
  assign link_sif_o_72_ = packet_i[17];
  assign link_sif_o[72] = link_sif_o_72_;
  assign link_sif_o_71_ = packet_i[16];
  assign link_sif_o[71] = link_sif_o_71_;
  assign link_sif_o_70_ = packet_i[15];
  assign link_sif_o[70] = link_sif_o_70_;
  assign link_sif_o_69_ = packet_i[14];
  assign link_sif_o[69] = link_sif_o_69_;
  assign link_sif_o_68_ = packet_i[13];
  assign link_sif_o[68] = link_sif_o_68_;
  assign link_sif_o_67_ = packet_i[12];
  assign link_sif_o[67] = link_sif_o_67_;
  assign link_sif_o_66_ = packet_i[11];
  assign link_sif_o[66] = link_sif_o_66_;
  assign link_sif_o_65_ = packet_i[10];
  assign link_sif_o[65] = link_sif_o_65_;
  assign link_sif_o_64_ = packet_i[9];
  assign link_sif_o[64] = link_sif_o_64_;
  assign link_sif_o_63_ = packet_i[8];
  assign link_sif_o[63] = link_sif_o_63_;
  assign link_sif_o_62_ = packet_i[7];
  assign link_sif_o[62] = link_sif_o_62_;
  assign link_sif_o_61_ = packet_i[6];
  assign link_sif_o[61] = link_sif_o_61_;
  assign link_sif_o_60_ = packet_i[5];
  assign link_sif_o[60] = link_sif_o_60_;
  assign link_sif_o_59_ = packet_i[4];
  assign link_sif_o[59] = link_sif_o_59_;
  assign link_sif_o_58_ = packet_i[3];
  assign link_sif_o[58] = link_sif_o_58_;
  assign link_sif_o_57_ = packet_i[2];
  assign link_sif_o[57] = link_sif_o_57_;
  assign link_sif_o_56_ = packet_i[1];
  assign link_sif_o[56] = link_sif_o_56_;
  assign link_sif_o_55_ = packet_i[0];
  assign link_sif_o[55] = link_sif_o_55_;
  assign link_sif_o_54_ = return_packet_v_i;
  assign link_sif_o[54] = link_sif_o_54_;
  assign link_sif_o_52_ = return_packet_i[52];
  assign link_sif_o[52] = link_sif_o_52_;
  assign link_sif_o_51_ = return_packet_i[51];
  assign link_sif_o[51] = link_sif_o_51_;
  assign link_sif_o_50_ = return_packet_i[50];
  assign link_sif_o[50] = link_sif_o_50_;
  assign link_sif_o_49_ = return_packet_i[49];
  assign link_sif_o[49] = link_sif_o_49_;
  assign link_sif_o_48_ = return_packet_i[48];
  assign link_sif_o[48] = link_sif_o_48_;
  assign link_sif_o_47_ = return_packet_i[47];
  assign link_sif_o[47] = link_sif_o_47_;
  assign link_sif_o_46_ = return_packet_i[46];
  assign link_sif_o[46] = link_sif_o_46_;
  assign link_sif_o_45_ = return_packet_i[45];
  assign link_sif_o[45] = link_sif_o_45_;
  assign link_sif_o_44_ = return_packet_i[44];
  assign link_sif_o[44] = link_sif_o_44_;
  assign link_sif_o_43_ = return_packet_i[43];
  assign link_sif_o[43] = link_sif_o_43_;
  assign link_sif_o_42_ = return_packet_i[42];
  assign link_sif_o[42] = link_sif_o_42_;
  assign link_sif_o_41_ = return_packet_i[41];
  assign link_sif_o[41] = link_sif_o_41_;
  assign link_sif_o_40_ = return_packet_i[40];
  assign link_sif_o[40] = link_sif_o_40_;
  assign link_sif_o_39_ = return_packet_i[39];
  assign link_sif_o[39] = link_sif_o_39_;
  assign link_sif_o_38_ = return_packet_i[38];
  assign link_sif_o[38] = link_sif_o_38_;
  assign link_sif_o_37_ = return_packet_i[37];
  assign link_sif_o[37] = link_sif_o_37_;
  assign link_sif_o_36_ = return_packet_i[36];
  assign link_sif_o[36] = link_sif_o_36_;
  assign link_sif_o_35_ = return_packet_i[35];
  assign link_sif_o[35] = link_sif_o_35_;
  assign link_sif_o_34_ = return_packet_i[34];
  assign link_sif_o[34] = link_sif_o_34_;
  assign link_sif_o_33_ = return_packet_i[33];
  assign link_sif_o[33] = link_sif_o_33_;
  assign link_sif_o_32_ = return_packet_i[32];
  assign link_sif_o[32] = link_sif_o_32_;
  assign link_sif_o_31_ = return_packet_i[31];
  assign link_sif_o[31] = link_sif_o_31_;
  assign link_sif_o_30_ = return_packet_i[30];
  assign link_sif_o[30] = link_sif_o_30_;
  assign link_sif_o_29_ = return_packet_i[29];
  assign link_sif_o[29] = link_sif_o_29_;
  assign link_sif_o_28_ = return_packet_i[28];
  assign link_sif_o[28] = link_sif_o_28_;
  assign link_sif_o_27_ = return_packet_i[27];
  assign link_sif_o[27] = link_sif_o_27_;
  assign link_sif_o_26_ = return_packet_i[26];
  assign link_sif_o[26] = link_sif_o_26_;
  assign link_sif_o_25_ = return_packet_i[25];
  assign link_sif_o[25] = link_sif_o_25_;
  assign link_sif_o_24_ = return_packet_i[24];
  assign link_sif_o[24] = link_sif_o_24_;
  assign link_sif_o_23_ = return_packet_i[23];
  assign link_sif_o[23] = link_sif_o_23_;
  assign link_sif_o_22_ = return_packet_i[22];
  assign link_sif_o[22] = link_sif_o_22_;
  assign link_sif_o_21_ = return_packet_i[21];
  assign link_sif_o[21] = link_sif_o_21_;
  assign link_sif_o_20_ = return_packet_i[20];
  assign link_sif_o[20] = link_sif_o_20_;
  assign link_sif_o_19_ = return_packet_i[19];
  assign link_sif_o[19] = link_sif_o_19_;
  assign link_sif_o_18_ = return_packet_i[18];
  assign link_sif_o[18] = link_sif_o_18_;
  assign link_sif_o_17_ = return_packet_i[17];
  assign link_sif_o[17] = link_sif_o_17_;
  assign link_sif_o_16_ = return_packet_i[16];
  assign link_sif_o[16] = link_sif_o_16_;
  assign link_sif_o_15_ = return_packet_i[15];
  assign link_sif_o[15] = link_sif_o_15_;
  assign link_sif_o_14_ = return_packet_i[14];
  assign link_sif_o[14] = link_sif_o_14_;
  assign link_sif_o_13_ = return_packet_i[13];
  assign link_sif_o[13] = link_sif_o_13_;
  assign link_sif_o_12_ = return_packet_i[12];
  assign link_sif_o[12] = link_sif_o_12_;
  assign link_sif_o_11_ = return_packet_i[11];
  assign link_sif_o[11] = link_sif_o_11_;
  assign link_sif_o_10_ = return_packet_i[10];
  assign link_sif_o[10] = link_sif_o_10_;
  assign link_sif_o_9_ = return_packet_i[9];
  assign link_sif_o[9] = link_sif_o_9_;
  assign link_sif_o_8_ = return_packet_i[8];
  assign link_sif_o[8] = link_sif_o_8_;
  assign link_sif_o_7_ = return_packet_i[7];
  assign link_sif_o[7] = link_sif_o_7_;
  assign link_sif_o_6_ = return_packet_i[6];
  assign link_sif_o[6] = link_sif_o_6_;
  assign link_sif_o_5_ = return_packet_i[5];
  assign link_sif_o[5] = link_sif_o_5_;
  assign link_sif_o_4_ = return_packet_i[4];
  assign link_sif_o[4] = link_sif_o_4_;
  assign link_sif_o_3_ = return_packet_i[3];
  assign link_sif_o[3] = link_sif_o_3_;
  assign link_sif_o_2_ = return_packet_i[2];
  assign link_sif_o[2] = link_sif_o_2_;
  assign link_sif_o_1_ = return_packet_i[1];
  assign link_sif_o[1] = link_sif_o_1_;
  assign link_sif_o_0_ = return_packet_i[0];
  assign link_sif_o[0] = link_sif_o_0_;

  bsg_fifo_1r1w_small_width_p97_els_p4
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(link_sif_i[153]),
    .ready_o(link_sif_o[152]),
    .data_i(link_sif_i[151:55]),
    .v_o(packet_v_o),
    .data_o(packet_o),
    .yumi_i(packet_yumi_i)
  );


  bsg_two_fifo_width_p53_allow_enq_deq_on_full_p1
  returned_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(returned_fifo_ready),
    .data_i(link_sif_i[52:0]),
    .v_i(link_sif_i[54]),
    .v_o(return_packet_v_o),
    .data_o(return_packet_o),
    .yumi_i(return_packet_yumi_i)
  );

  assign return_packet_fifo_full_o = ~returned_fifo_ready;

endmodule



module bsg_counter_up_down_max_val_p63_init_val_p0_max_step_p1
(
  clk_i,
  reset_i,
  up_i,
  down_i,
  count_o
);

  input [0:0] up_i;
  input [0:0] down_i;
  output [5:0] count_o;
  input clk_i;
  input reset_i;
  wire [5:0] count_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;
  reg count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,count_o_2_sv2v_reg,
  count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign { N6, N5, N4, N3, N2, N1 } = count_o - down_i[0];
  assign { N12, N11, N10, N9, N8, N7 } = { N6, N5, N4, N3, N2, N1 } + up_i[0];
  assign N0 = ~reset_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
      count_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_5_sv2v_reg <= N12;
      count_o_4_sv2v_reg <= N11;
      count_o_3_sv2v_reg <= N10;
      count_o_2_sv2v_reg <= N9;
      count_o_1_sv2v_reg <= N8;
      count_o_0_sv2v_reg <= N7;
    end 
  end


endmodule



module bsg_manycore_endpoint_fc_x_cord_width_p7_y_cord_width_p7_fifo_els_p4_data_width_p32_addr_width_p28_credit_counter_width_p6_warn_out_of_credits_p1_rev_fifo_els_p2_use_credits_for_local_fifo_p1
(
  clk_i,
  reset_i,
  link_sif_i,
  link_sif_o,
  packet_o,
  packet_v_o,
  packet_yumi_i,
  return_packet_i,
  return_packet_v_i,
  packet_i,
  packet_v_i,
  packet_credit_or_ready_o,
  return_packet_o,
  return_packet_v_o,
  return_packet_yumi_i,
  return_packet_fifo_full_o,
  out_credits_used_o
);

  input [153:0] link_sif_i;
  output [153:0] link_sif_o;
  output [96:0] packet_o;
  input [52:0] return_packet_i;
  input [96:0] packet_i;
  output [52:0] return_packet_o;
  output [5:0] out_credits_used_o;
  input clk_i;
  input reset_i;
  input packet_yumi_i;
  input return_packet_v_i;
  input packet_v_i;
  input return_packet_yumi_i;
  output packet_v_o;
  output packet_credit_or_ready_o;
  output return_packet_v_o;
  output return_packet_fifo_full_o;
  wire [153:0] link_sif_o;
  wire [96:0] packet_o;
  wire [52:0] return_packet_o;
  wire [5:0] out_credits_used_o;
  wire packet_v_o,packet_credit_or_ready_o,return_packet_v_o,return_packet_fifo_full_o,
  packet_v_lo,return_packet_credit_or_ready_lo,rev_fifo_has_space,N0,N1,N2,N3,
  returned_credit;
  wire [1:0] rev_fifo_credit_r,rev_fifo_credit_available;
  reg rev_fifo_credit_r_1_sv2v_reg,rev_fifo_credit_r_0_sv2v_reg;
  assign rev_fifo_credit_r[1] = rev_fifo_credit_r_1_sv2v_reg;
  assign rev_fifo_credit_r[0] = rev_fifo_credit_r_0_sv2v_reg;

  bsg_manycore_endpoint_x_cord_width_p7_y_cord_width_p7_fifo_els_p4_data_width_p32_addr_width_p28
  bme
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_sif_i(link_sif_i),
    .link_sif_o(link_sif_o),
    .packet_o(packet_o),
    .packet_v_o(packet_v_lo),
    .packet_yumi_i(packet_yumi_i),
    .return_packet_i(return_packet_i),
    .return_packet_v_i(return_packet_v_i),
    .return_packet_credit_or_ready_o(return_packet_credit_or_ready_lo),
    .packet_i(packet_i),
    .packet_v_i(packet_v_i),
    .packet_credit_or_ready_o(packet_credit_or_ready_o),
    .return_packet_o(return_packet_o),
    .return_packet_v_o(return_packet_v_o),
    .return_packet_yumi_i(return_packet_yumi_i),
    .return_packet_fifo_full_o(return_packet_fifo_full_o)
  );

  assign rev_fifo_has_space = rev_fifo_credit_available != 1'b0;

  bsg_counter_up_down_max_val_p63_init_val_p0_max_step_p1
  out_credit_ctr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .up_i(packet_v_i),
    .down_i(returned_credit),
    .count_o(out_credits_used_o)
  );

  assign rev_fifo_credit_available = rev_fifo_credit_r + return_packet_credit_or_ready_lo;
  assign { N3, N2 } = rev_fifo_credit_available - N1;
  assign N0 = ~reset_i;
  assign N1 = packet_v_lo & packet_yumi_i;
  assign packet_v_o = packet_v_lo & rev_fifo_has_space;
  assign returned_credit = return_packet_v_o & return_packet_yumi_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      rev_fifo_credit_r_1_sv2v_reg <= 1'b1;
      rev_fifo_credit_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      rev_fifo_credit_r_1_sv2v_reg <= N3;
      rev_fifo_credit_r_0_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_manycore_reg_id_decode
(
  data_i,
  mask_i,
  reg_id_o
);

  input [31:0] data_i;
  input [3:0] mask_i;
  output [4:0] reg_id_o;
  wire [4:0] reg_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33;
  assign reg_id_o[4] = N7 | N9;
  assign N7 = N4 | N6;
  assign N4 = N1 | N3;
  assign N1 = data_i[4] & N0;
  assign N0 = ~mask_i[0];
  assign N3 = data_i[12] & N2;
  assign N2 = ~mask_i[1];
  assign N6 = data_i[20] & N5;
  assign N5 = ~mask_i[2];
  assign N9 = data_i[28] & N8;
  assign N8 = ~mask_i[3];
  assign reg_id_o[3] = N14 | N15;
  assign N14 = N12 | N13;
  assign N12 = N10 | N11;
  assign N10 = data_i[3] & N0;
  assign N11 = data_i[11] & N2;
  assign N13 = data_i[19] & N5;
  assign N15 = data_i[27] & N8;
  assign reg_id_o[2] = N20 | N21;
  assign N20 = N18 | N19;
  assign N18 = N16 | N17;
  assign N16 = data_i[2] & N0;
  assign N17 = data_i[10] & N2;
  assign N19 = data_i[18] & N5;
  assign N21 = data_i[26] & N8;
  assign reg_id_o[1] = N26 | N27;
  assign N26 = N24 | N25;
  assign N24 = N22 | N23;
  assign N22 = data_i[1] & N0;
  assign N23 = data_i[9] & N2;
  assign N25 = data_i[17] & N5;
  assign N27 = data_i[25] & N8;
  assign reg_id_o[0] = N32 | N33;
  assign N32 = N30 | N31;
  assign N30 = N28 | N29;
  assign N28 = data_i[0] & N0;
  assign N29 = data_i[8] & N2;
  assign N31 = data_i[16] & N5;
  assign N33 = data_i[24] & N8;

endmodule



module bsg_manycore_endpoint_standard_x_cord_width_p7_y_cord_width_p7_fifo_els_p4_data_width_p32_addr_width_p28_credit_counter_width_p6_rev_fifo_els_p2_use_credits_for_local_fifo_p1
(
  clk_i,
  reset_i,
  link_sif_i,
  link_sif_o,
  in_v_o,
  in_data_o,
  in_mask_o,
  in_addr_o,
  in_we_o,
  in_load_info_o,
  in_src_x_cord_o,
  in_src_y_cord_o,
  in_yumi_i,
  returning_data_i,
  returning_v_i,
  out_v_i,
  out_packet_i,
  out_credit_or_ready_o,
  returned_data_r_o,
  returned_reg_id_r_o,
  returned_v_r_o,
  returned_pkt_type_r_o,
  returned_yumi_i,
  returned_fifo_full_o,
  returned_credit_v_r_o,
  returned_credit_reg_id_r_o,
  out_credits_used_o,
  global_x_i,
  global_y_i
);

  input [153:0] link_sif_i;
  output [153:0] link_sif_o;
  output [31:0] in_data_o;
  output [3:0] in_mask_o;
  output [27:0] in_addr_o;
  output [6:0] in_load_info_o;
  output [6:0] in_src_x_cord_o;
  output [6:0] in_src_y_cord_o;
  input [31:0] returning_data_i;
  input [96:0] out_packet_i;
  output [31:0] returned_data_r_o;
  output [4:0] returned_reg_id_r_o;
  output [1:0] returned_pkt_type_r_o;
  output [4:0] returned_credit_reg_id_r_o;
  output [5:0] out_credits_used_o;
  input [6:0] global_x_i;
  input [6:0] global_y_i;
  input clk_i;
  input reset_i;
  input in_yumi_i;
  input returning_v_i;
  input out_v_i;
  input returned_yumi_i;
  output in_v_o;
  output in_we_o;
  output out_credit_or_ready_o;
  output returned_v_r_o;
  output returned_fifo_full_o;
  output returned_credit_v_r_o;
  wire [153:0] link_sif_o;
  wire [31:0] in_data_o,returned_data_r_o;
  wire [3:0] in_mask_o;
  wire [27:0] in_addr_o;
  wire [6:0] in_load_info_o,in_src_x_cord_o,in_src_y_cord_o;
  wire [4:0] returned_reg_id_r_o,returned_credit_reg_id_r_o,payload_reg_id,return_reg_id;
  wire [1:0] returned_pkt_type_r_o,return_pkt_type;
  wire [5:0] out_credits_used_o;
  wire in_v_o,in_we_o,out_credit_or_ready_o,returned_v_r_o,returned_fifo_full_o,
  returned_credit_v_r_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,in_data_o_6_,in_data_o_5_,
  in_data_o_4_,in_data_o_3_,in_data_o_2_,in_data_o_1_,in_data_o_0_,packet_lo_op_v2__3_,
  packet_lo_op_v2__2_,packet_lo_op_v2__1_,packet_lo_op_v2__0_,packet_lo_reg_id__4_,
  packet_lo_reg_id__3_,packet_lo_reg_id__2_,packet_lo_reg_id__1_,packet_lo_reg_id__0_,
  packet_lo_y_cord__6_,packet_lo_y_cord__5_,packet_lo_y_cord__4_,
  packet_lo_y_cord__3_,packet_lo_y_cord__2_,packet_lo_y_cord__1_,packet_lo_y_cord__0_,
  packet_lo_x_cord__6_,packet_lo_x_cord__5_,packet_lo_x_cord__4_,packet_lo_x_cord__3_,
  packet_lo_x_cord__2_,packet_lo_x_cord__1_,packet_lo_x_cord__0_,packet_v_lo,packet_yumi_li,
  return_packet_li_data__31_,return_packet_li_data__30_,return_packet_li_data__29_,
  return_packet_li_data__28_,return_packet_li_data__27_,
  return_packet_li_data__26_,return_packet_li_data__25_,return_packet_li_data__24_,
  return_packet_li_data__23_,return_packet_li_data__22_,return_packet_li_data__21_,
  return_packet_li_data__20_,return_packet_li_data__19_,return_packet_li_data__18_,
  return_packet_li_data__17_,return_packet_li_data__16_,return_packet_li_data__15_,
  return_packet_li_data__14_,return_packet_li_data__13_,return_packet_li_data__12_,
  return_packet_li_data__11_,return_packet_li_data__10_,return_packet_li_data__9_,
  return_packet_li_data__8_,return_packet_li_data__7_,return_packet_li_data__6_,
  return_packet_li_data__5_,return_packet_li_data__4_,return_packet_li_data__3_,
  return_packet_li_data__2_,return_packet_li_data__1_,return_packet_li_data__0_,return_packet_v_li,
  return_packet_lo_y_cord__6_,return_packet_lo_y_cord__5_,return_packet_lo_y_cord__4_,
  return_packet_lo_y_cord__3_,return_packet_lo_y_cord__2_,return_packet_lo_y_cord__1_,
  return_packet_lo_y_cord__0_,return_packet_lo_x_cord__6_,
  return_packet_lo_x_cord__5_,return_packet_lo_x_cord__4_,return_packet_lo_x_cord__3_,
  return_packet_lo_x_cord__2_,return_packet_lo_x_cord__1_,return_packet_lo_x_cord__0_,
  return_packet_v_lo,return_packet_yumi_li,lock_r,lock_v_r,lock_return_r,lock_n,lock_v_n,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,
  N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46;
  wire [20:0] return_info_r;
  reg lock_return_r_sv2v_reg,lock_r_sv2v_reg,lock_v_r_sv2v_reg,
  return_info_r_20_sv2v_reg,return_info_r_19_sv2v_reg,return_info_r_18_sv2v_reg,
  return_info_r_17_sv2v_reg,return_info_r_16_sv2v_reg,return_info_r_15_sv2v_reg,return_info_r_14_sv2v_reg,
  return_info_r_13_sv2v_reg,return_info_r_12_sv2v_reg,return_info_r_11_sv2v_reg,
  return_info_r_10_sv2v_reg,return_info_r_9_sv2v_reg,return_info_r_8_sv2v_reg,
  return_info_r_7_sv2v_reg,return_info_r_6_sv2v_reg,return_info_r_5_sv2v_reg,
  return_info_r_4_sv2v_reg,return_info_r_3_sv2v_reg,return_info_r_2_sv2v_reg,
  return_info_r_1_sv2v_reg,return_info_r_0_sv2v_reg;
  assign lock_return_r = lock_return_r_sv2v_reg;
  assign lock_r = lock_r_sv2v_reg;
  assign lock_v_r = lock_v_r_sv2v_reg;
  assign return_info_r[20] = return_info_r_20_sv2v_reg;
  assign return_info_r[19] = return_info_r_19_sv2v_reg;
  assign return_info_r[18] = return_info_r_18_sv2v_reg;
  assign return_info_r[17] = return_info_r_17_sv2v_reg;
  assign return_info_r[16] = return_info_r_16_sv2v_reg;
  assign return_info_r[15] = return_info_r_15_sv2v_reg;
  assign return_info_r[14] = return_info_r_14_sv2v_reg;
  assign return_info_r[13] = return_info_r_13_sv2v_reg;
  assign return_info_r[12] = return_info_r_12_sv2v_reg;
  assign return_info_r[11] = return_info_r_11_sv2v_reg;
  assign return_info_r[10] = return_info_r_10_sv2v_reg;
  assign return_info_r[9] = return_info_r_9_sv2v_reg;
  assign return_info_r[8] = return_info_r_8_sv2v_reg;
  assign return_info_r[7] = return_info_r_7_sv2v_reg;
  assign return_info_r[6] = return_info_r_6_sv2v_reg;
  assign return_info_r[5] = return_info_r_5_sv2v_reg;
  assign return_info_r[4] = return_info_r_4_sv2v_reg;
  assign return_info_r[3] = return_info_r_3_sv2v_reg;
  assign return_info_r[2] = return_info_r_2_sv2v_reg;
  assign return_info_r[1] = return_info_r_1_sv2v_reg;
  assign return_info_r[0] = return_info_r_0_sv2v_reg;
  assign in_load_info_o[6] = in_data_o_6_;
  assign in_data_o[6] = in_data_o_6_;
  assign in_load_info_o[5] = in_data_o_5_;
  assign in_data_o[5] = in_data_o_5_;
  assign in_load_info_o[4] = in_data_o_4_;
  assign in_data_o[4] = in_data_o_4_;
  assign in_load_info_o[3] = in_data_o_3_;
  assign in_data_o[3] = in_data_o_3_;
  assign in_load_info_o[2] = in_data_o_2_;
  assign in_data_o[2] = in_data_o_2_;
  assign in_load_info_o[1] = in_data_o_1_;
  assign in_data_o[1] = in_data_o_1_;
  assign in_load_info_o[0] = in_data_o_0_;
  assign in_data_o[0] = in_data_o_0_;
  assign returned_credit_reg_id_r_o[4] = returned_reg_id_r_o[4];
  assign returned_credit_reg_id_r_o[3] = returned_reg_id_r_o[3];
  assign returned_credit_reg_id_r_o[2] = returned_reg_id_r_o[2];
  assign returned_credit_reg_id_r_o[1] = returned_reg_id_r_o[1];
  assign returned_credit_reg_id_r_o[0] = returned_reg_id_r_o[0];

  bsg_manycore_endpoint_fc_x_cord_width_p7_y_cord_width_p7_fifo_els_p4_data_width_p32_addr_width_p28_credit_counter_width_p6_warn_out_of_credits_p1_rev_fifo_els_p2_use_credits_for_local_fifo_p1
  bme
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_sif_i(link_sif_i),
    .link_sif_o(link_sif_o),
    .packet_o({ in_addr_o, packet_lo_op_v2__3_, packet_lo_op_v2__2_, packet_lo_op_v2__1_, packet_lo_op_v2__0_, packet_lo_reg_id__4_, packet_lo_reg_id__3_, packet_lo_reg_id__2_, packet_lo_reg_id__1_, packet_lo_reg_id__0_, in_data_o[31:7], in_data_o_6_, in_data_o_5_, in_data_o_4_, in_data_o_3_, in_data_o_2_, in_data_o_1_, in_data_o_0_, in_src_y_cord_o, in_src_x_cord_o, packet_lo_y_cord__6_, packet_lo_y_cord__5_, packet_lo_y_cord__4_, packet_lo_y_cord__3_, packet_lo_y_cord__2_, packet_lo_y_cord__1_, packet_lo_y_cord__0_, packet_lo_x_cord__6_, packet_lo_x_cord__5_, packet_lo_x_cord__4_, packet_lo_x_cord__3_, packet_lo_x_cord__2_, packet_lo_x_cord__1_, packet_lo_x_cord__0_ }),
    .packet_v_o(packet_v_lo),
    .packet_yumi_i(packet_yumi_li),
    .return_packet_i({ return_info_r[1:0], return_packet_li_data__31_, return_packet_li_data__30_, return_packet_li_data__29_, return_packet_li_data__28_, return_packet_li_data__27_, return_packet_li_data__26_, return_packet_li_data__25_, return_packet_li_data__24_, return_packet_li_data__23_, return_packet_li_data__22_, return_packet_li_data__21_, return_packet_li_data__20_, return_packet_li_data__19_, return_packet_li_data__18_, return_packet_li_data__17_, return_packet_li_data__16_, return_packet_li_data__15_, return_packet_li_data__14_, return_packet_li_data__13_, return_packet_li_data__12_, return_packet_li_data__11_, return_packet_li_data__10_, return_packet_li_data__9_, return_packet_li_data__8_, return_packet_li_data__7_, return_packet_li_data__6_, return_packet_li_data__5_, return_packet_li_data__4_, return_packet_li_data__3_, return_packet_li_data__2_, return_packet_li_data__1_, return_packet_li_data__0_, return_info_r[6:2], return_info_r[20:7] }),
    .return_packet_v_i(return_packet_v_li),
    .packet_i(out_packet_i),
    .packet_v_i(out_v_i),
    .packet_credit_or_ready_o(out_credit_or_ready_o),
    .return_packet_o({ returned_pkt_type_r_o, returned_data_r_o, returned_reg_id_r_o, return_packet_lo_y_cord__6_, return_packet_lo_y_cord__5_, return_packet_lo_y_cord__4_, return_packet_lo_y_cord__3_, return_packet_lo_y_cord__2_, return_packet_lo_y_cord__1_, return_packet_lo_y_cord__0_, return_packet_lo_x_cord__6_, return_packet_lo_x_cord__5_, return_packet_lo_x_cord__4_, return_packet_lo_x_cord__3_, return_packet_lo_x_cord__2_, return_packet_lo_x_cord__1_, return_packet_lo_x_cord__0_ }),
    .return_packet_v_o(return_packet_v_lo),
    .return_packet_yumi_i(return_packet_yumi_li),
    .return_packet_fifo_full_o(returned_fifo_full_o),
    .out_credits_used_o(out_credits_used_o)
  );


  bsg_manycore_reg_id_decode
  pd0
  (
    .data_i({ in_data_o[31:7], in_data_o_6_, in_data_o_5_, in_data_o_4_, in_data_o_3_, in_data_o_2_, in_data_o_1_, in_data_o_0_ }),
    .mask_i({ packet_lo_reg_id__3_, packet_lo_reg_id__2_, packet_lo_reg_id__1_, packet_lo_reg_id__0_ }),
    .reg_id_o(payload_reg_id)
  );

  assign N13 = N9 & N10;
  assign N14 = N11 & N12;
  assign N15 = N13 & N14;
  assign N16 = packet_lo_op_v2__3_ | packet_lo_op_v2__2_;
  assign N17 = N11 | packet_lo_op_v2__0_;
  assign N18 = N16 | N17;
  assign N20 = packet_lo_op_v2__3_ | packet_lo_op_v2__2_;
  assign N21 = packet_lo_op_v2__1_ | N12;
  assign N22 = N20 | N21;
  assign N24 = packet_lo_op_v2__3_ | N10;
  assign N25 = packet_lo_op_v2__1_ | packet_lo_op_v2__0_;
  assign N26 = N24 | N25;
  assign N28 = packet_lo_op_v2__2_ & packet_lo_op_v2__0_;
  assign N29 = packet_lo_op_v2__1_ & packet_lo_op_v2__0_;
  assign N30 = packet_lo_op_v2__2_ & packet_lo_op_v2__1_;
  assign N40 = reset_i | N15;
  assign N41 = returned_pkt_type_r_o[0] | returned_pkt_type_r_o[1];
  assign N42 = returned_pkt_type_r_o[0] | returned_pkt_type_r_o[1];
  assign N43 = ~N42;
  assign N32 = ~N33;
  assign N35 = (N0)? in_data_o_0_ : 
               (N1)? lock_r : 1'b0;
  assign N0 = packet_v_lo;
  assign N1 = N34;
  assign in_v_o = (N2)? packet_v_lo : 
                  (N3)? packet_v_lo : 
                  (N4)? packet_v_lo : 
                  (N5)? 1'b0 : 
                  (N6)? 1'b0 : 1'b0;
  assign N2 = N15;
  assign N3 = N19;
  assign N4 = N23;
  assign N5 = N27;
  assign N6 = N31;
  assign packet_yumi_li = (N2)? in_yumi_i : 
                          (N3)? in_yumi_i : 
                          (N4)? in_yumi_i : 
                          (N5)? packet_v_lo : 
                          (N6)? 1'b0 : 1'b0;
  assign return_pkt_type[0] = (N2)? N32 : 
                              (N3)? 1'b0 : 
                              (N4)? 1'b0 : 
                              (N5)? 1'b1 : 
                              (N6)? 1'b0 : 1'b0;
  assign return_pkt_type[1] = (N2)? N33 : 
                              (N37)? 1'b0 : 1'b0;
  assign in_we_o = (N2)? 1'b0 : 
                   (N3)? 1'b1 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b0 : 
                   (N6)? 1'b0 : 1'b0;
  assign in_mask_o = (N2)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                     (N3)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                     (N4)? { packet_lo_reg_id__3_, packet_lo_reg_id__2_, packet_lo_reg_id__1_, packet_lo_reg_id__0_ } : 
                     (N5)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                     (N6)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign return_reg_id = (N2)? { packet_lo_reg_id__4_, packet_lo_reg_id__3_, packet_lo_reg_id__2_, packet_lo_reg_id__1_, packet_lo_reg_id__0_ } : 
                         (N3)? { packet_lo_reg_id__4_, packet_lo_reg_id__3_, packet_lo_reg_id__2_, packet_lo_reg_id__1_, packet_lo_reg_id__0_ } : 
                         (N4)? payload_reg_id : 
                         (N5)? { packet_lo_reg_id__4_, packet_lo_reg_id__3_, packet_lo_reg_id__2_, packet_lo_reg_id__1_, packet_lo_reg_id__0_ } : 
                         (N6)? { packet_lo_reg_id__4_, packet_lo_reg_id__3_, packet_lo_reg_id__2_, packet_lo_reg_id__1_, packet_lo_reg_id__0_ } : 1'b0;
  assign lock_v_n = (N3)? 1'b0 : 
                    (N4)? 1'b0 : 
                    (N5)? packet_v_lo : 
                    (N6)? 1'b0 : 1'b0;
  assign lock_n = (N2)? lock_r : 
                  (N3)? lock_r : 
                  (N4)? lock_r : 
                  (N5)? N35 : 
                  (N6)? lock_r : 1'b0;
  assign { return_packet_li_data__31_, return_packet_li_data__30_, return_packet_li_data__29_, return_packet_li_data__28_, return_packet_li_data__27_, return_packet_li_data__26_, return_packet_li_data__25_, return_packet_li_data__24_, return_packet_li_data__23_, return_packet_li_data__22_, return_packet_li_data__21_, return_packet_li_data__20_, return_packet_li_data__19_, return_packet_li_data__18_, return_packet_li_data__17_, return_packet_li_data__16_, return_packet_li_data__15_, return_packet_li_data__14_, return_packet_li_data__13_, return_packet_li_data__12_, return_packet_li_data__11_, return_packet_li_data__10_, return_packet_li_data__9_, return_packet_li_data__8_, return_packet_li_data__7_, return_packet_li_data__6_, return_packet_li_data__5_, return_packet_li_data__4_, return_packet_li_data__3_, return_packet_li_data__2_, return_packet_li_data__1_, return_packet_li_data__0_ } = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lock_return_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N8)? returning_data_i : 1'b0;
  assign N7 = lock_v_r;
  assign N8 = N39;
  assign N9 = ~packet_lo_op_v2__3_;
  assign N10 = ~packet_lo_op_v2__2_;
  assign N11 = ~packet_lo_op_v2__1_;
  assign N12 = ~packet_lo_op_v2__0_;
  assign N19 = ~N18;
  assign N23 = ~N22;
  assign N27 = ~N26;
  assign N31 = packet_lo_op_v2__3_ | N45;
  assign N45 = N28 | N44;
  assign N44 = N29 | N30;
  assign N33 = in_data_o_6_;
  assign N34 = ~packet_v_lo;
  assign N36 = ~N15;
  assign N37 = N36;
  assign N38 = packet_v_lo & packet_yumi_li;
  assign return_packet_v_li = lock_v_r | returning_v_i;
  assign N39 = ~lock_v_r;
  assign returned_v_r_o = return_packet_v_lo & N41;
  assign return_packet_yumi_li = returned_yumi_i | N46;
  assign N46 = return_packet_v_lo & N43;
  assign returned_credit_v_r_o = return_packet_v_lo & return_packet_yumi_li;

  always @(posedge clk_i) begin
    if(reset_i) begin
      lock_return_r_sv2v_reg <= 1'b0;
      lock_r_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      lock_return_r_sv2v_reg <= lock_r;
      lock_r_sv2v_reg <= lock_n;
    end 
    if(N40) begin
      lock_v_r_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      lock_v_r_sv2v_reg <= lock_v_n;
    end 
    if(N38) begin
      return_info_r_20_sv2v_reg <= in_src_y_cord_o[6];
      return_info_r_19_sv2v_reg <= in_src_y_cord_o[5];
      return_info_r_18_sv2v_reg <= in_src_y_cord_o[4];
      return_info_r_17_sv2v_reg <= in_src_y_cord_o[3];
      return_info_r_16_sv2v_reg <= in_src_y_cord_o[2];
      return_info_r_15_sv2v_reg <= in_src_y_cord_o[1];
      return_info_r_14_sv2v_reg <= in_src_y_cord_o[0];
      return_info_r_13_sv2v_reg <= in_src_x_cord_o[6];
      return_info_r_12_sv2v_reg <= in_src_x_cord_o[5];
      return_info_r_11_sv2v_reg <= in_src_x_cord_o[4];
      return_info_r_10_sv2v_reg <= in_src_x_cord_o[3];
      return_info_r_9_sv2v_reg <= in_src_x_cord_o[2];
      return_info_r_8_sv2v_reg <= in_src_x_cord_o[1];
      return_info_r_7_sv2v_reg <= in_src_x_cord_o[0];
      return_info_r_6_sv2v_reg <= return_reg_id[4];
      return_info_r_5_sv2v_reg <= return_reg_id[3];
      return_info_r_4_sv2v_reg <= return_reg_id[2];
      return_info_r_3_sv2v_reg <= return_reg_id[1];
      return_info_r_2_sv2v_reg <= return_reg_id[0];
      return_info_r_1_sv2v_reg <= return_pkt_type[1];
      return_info_r_0_sv2v_reg <= return_pkt_type[0];
    end 
  end


endmodule



module bsg_mux_width_p8_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [1:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[15] : 
                     (N3)? data_i[23] : 
                     (N5)? data_i[31] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[14] : 
                     (N3)? data_i[22] : 
                     (N5)? data_i[30] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[13] : 
                     (N3)? data_i[21] : 
                     (N5)? data_i[29] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[12] : 
                     (N3)? data_i[20] : 
                     (N5)? data_i[28] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[11] : 
                     (N3)? data_i[19] : 
                     (N5)? data_i[27] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[10] : 
                     (N3)? data_i[18] : 
                     (N5)? data_i[26] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[9] : 
                     (N3)? data_i[17] : 
                     (N5)? data_i[25] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[8] : 
                     (N3)? data_i[16] : 
                     (N5)? data_i[24] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p16_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [0:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[31] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[30] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[29] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[28] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[27] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[26] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[25] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[24] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[23] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[22] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[21] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[20] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[19] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[18] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[17] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[16] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module load_packer
(
  mem_data_i,
  unsigned_load_i,
  byte_load_i,
  hex_load_i,
  part_sel_i,
  load_data_o
);

  input [31:0] mem_data_i;
  input [1:0] part_sel_i;
  output [31:0] load_data_o;
  input unsigned_load_i;
  input byte_load_i;
  input hex_load_i;
  wire [31:0] load_data_o;
  wire N0,half_sigext,byte_sigext,N1,N2,N3,N4,N5;
  wire [7:0] loaded_byte;
  wire [15:0] loaded_half;

  bsg_mux_width_p8_els_p4
  byte_sel_mux
  (
    .data_i(mem_data_i),
    .sel_i(part_sel_i),
    .data_o(loaded_byte)
  );


  bsg_mux_width_p16_els_p2
  half_sel_mux
  (
    .data_i(mem_data_i),
    .sel_i(part_sel_i[1]),
    .data_o(loaded_half)
  );

  assign load_data_o = (N0)? { byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, byte_sigext, loaded_byte } : 
                       (N4)? { half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, half_sigext, loaded_half } : 
                       (N2)? mem_data_i : 1'b0;
  assign N0 = byte_load_i;
  assign half_sigext = N5 & loaded_half[15];
  assign N5 = ~unsigned_load_i;
  assign byte_sigext = N5 & loaded_byte[7];
  assign N1 = hex_load_i | byte_load_i;
  assign N2 = ~N1;
  assign N3 = ~byte_load_i;
  assign N4 = hex_load_i & N3;

endmodule



module network_rx_data_width_p32_addr_width_p28_dmem_size_p1024_icache_tag_width_p12_icache_entries_p1024_x_cord_width_p7_y_cord_width_p7_x_subcord_width_p4_y_subcord_width_p3
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  mask_i,
  load_info_i,
  yumi_o,
  src_x_cord_debug_i,
  src_y_cord_debug_i,
  returning_data_o,
  returning_data_v_o,
  remote_dmem_v_o,
  remote_dmem_w_o,
  remote_dmem_addr_o,
  remote_dmem_mask_o,
  remote_dmem_data_o,
  remote_dmem_data_i,
  remote_dmem_yumi_i,
  icache_v_o,
  icache_pc_o,
  icache_instr_o,
  icache_yumi_i,
  freeze_o,
  tgo_x_o,
  tgo_y_o,
  pc_init_val_o,
  remote_interrupt_set_o,
  remote_interrupt_clear_o,
  remote_interrupt_pending_bit_i,
  global_x_i,
  global_y_i
);

  input [27:0] addr_i;
  input [31:0] data_i;
  input [3:0] mask_i;
  input [6:0] load_info_i;
  input [6:0] src_x_cord_debug_i;
  input [6:0] src_y_cord_debug_i;
  output [31:0] returning_data_o;
  output [9:0] remote_dmem_addr_o;
  output [3:0] remote_dmem_mask_o;
  output [31:0] remote_dmem_data_o;
  input [31:0] remote_dmem_data_i;
  output [21:0] icache_pc_o;
  output [31:0] icache_instr_o;
  output [3:0] tgo_x_o;
  output [2:0] tgo_y_o;
  output [21:0] pc_init_val_o;
  input [6:0] global_x_i;
  input [6:0] global_y_i;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  input remote_dmem_yumi_i;
  input icache_yumi_i;
  input remote_interrupt_pending_bit_i;
  output yumi_o;
  output returning_data_v_o;
  output remote_dmem_v_o;
  output remote_dmem_w_o;
  output icache_v_o;
  output freeze_o;
  output remote_interrupt_set_o;
  output remote_interrupt_clear_o;
  wire [31:0] returning_data_o,remote_dmem_data_o,icache_instr_o,load_data_lo;
  wire [9:0] remote_dmem_addr_o;
  wire [3:0] remote_dmem_mask_o,tgo_x_o;
  wire [21:0] icache_pc_o,pc_init_val_o;
  wire [2:0] tgo_y_o;
  wire yumi_o,returning_data_v_o,remote_dmem_v_o,remote_dmem_w_o,icache_v_o,freeze_o,
  remote_interrupt_set_o,remote_interrupt_clear_o,N0,N1,N2,N3,N4,N5,N6,
  icache_pc_o_21_,icache_pc_o_20_,icache_pc_o_19_,icache_pc_o_18_,icache_pc_o_17_,
  icache_pc_o_16_,icache_pc_o_15_,icache_pc_o_14_,icache_pc_o_13_,icache_pc_o_12_,
  icache_pc_o_11_,icache_pc_o_10_,is_icache_addr,is_csr_addr,is_freeze_addr,is_tgo_x_addr,
  is_tgo_y_addr,is_pc_init_val_addr,load_info_r_is_unsigned_op_,
  load_info_r_is_byte_op_,load_info_r_is_hex_op_,load_info_r_part_sel__1_,load_info_r_part_sel__0_,N7,N8,
  N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,
  N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,
  N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,
  N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,
  N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,
  N107,send_dmem_data_r,send_freeze_r,send_tgo_x_r,send_tgo_y_r,send_pc_init_val_r,
  send_invalid_r,send_zero_r,send_remote_interrupt_r,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,
  N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
  N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,
  N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,
  N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,
  N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,
  N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,
  N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
  N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,
  N306,N307,N308,N309,N310;
  reg load_info_r_is_unsigned_op__sv2v_reg,load_info_r_is_byte_op__sv2v_reg,
  load_info_r_is_hex_op__sv2v_reg,load_info_r_part_sel__1__sv2v_reg,
  load_info_r_part_sel__0__sv2v_reg,freeze_o_sv2v_reg,tgo_x_o_3_sv2v_reg,tgo_x_o_2_sv2v_reg,
  tgo_x_o_1_sv2v_reg,tgo_x_o_0_sv2v_reg,tgo_y_o_2_sv2v_reg,tgo_y_o_1_sv2v_reg,
  tgo_y_o_0_sv2v_reg,pc_init_val_o_21_sv2v_reg,pc_init_val_o_20_sv2v_reg,pc_init_val_o_19_sv2v_reg,
  pc_init_val_o_18_sv2v_reg,pc_init_val_o_17_sv2v_reg,pc_init_val_o_16_sv2v_reg,
  pc_init_val_o_15_sv2v_reg,pc_init_val_o_14_sv2v_reg,pc_init_val_o_13_sv2v_reg,
  pc_init_val_o_12_sv2v_reg,pc_init_val_o_11_sv2v_reg,pc_init_val_o_10_sv2v_reg,
  pc_init_val_o_9_sv2v_reg,pc_init_val_o_8_sv2v_reg,pc_init_val_o_7_sv2v_reg,
  pc_init_val_o_6_sv2v_reg,pc_init_val_o_5_sv2v_reg,pc_init_val_o_4_sv2v_reg,
  pc_init_val_o_3_sv2v_reg,pc_init_val_o_2_sv2v_reg,pc_init_val_o_1_sv2v_reg,
  pc_init_val_o_0_sv2v_reg,send_dmem_data_r_sv2v_reg,send_freeze_r_sv2v_reg,send_tgo_x_r_sv2v_reg,
  send_tgo_y_r_sv2v_reg,send_pc_init_val_r_sv2v_reg,send_invalid_r_sv2v_reg,
  send_zero_r_sv2v_reg,send_remote_interrupt_r_sv2v_reg;
  assign load_info_r_is_unsigned_op_ = load_info_r_is_unsigned_op__sv2v_reg;
  assign load_info_r_is_byte_op_ = load_info_r_is_byte_op__sv2v_reg;
  assign load_info_r_is_hex_op_ = load_info_r_is_hex_op__sv2v_reg;
  assign load_info_r_part_sel__1_ = load_info_r_part_sel__1__sv2v_reg;
  assign load_info_r_part_sel__0_ = load_info_r_part_sel__0__sv2v_reg;
  assign freeze_o = freeze_o_sv2v_reg;
  assign tgo_x_o[3] = tgo_x_o_3_sv2v_reg;
  assign tgo_x_o[2] = tgo_x_o_2_sv2v_reg;
  assign tgo_x_o[1] = tgo_x_o_1_sv2v_reg;
  assign tgo_x_o[0] = tgo_x_o_0_sv2v_reg;
  assign tgo_y_o[2] = tgo_y_o_2_sv2v_reg;
  assign tgo_y_o[1] = tgo_y_o_1_sv2v_reg;
  assign tgo_y_o[0] = tgo_y_o_0_sv2v_reg;
  assign pc_init_val_o[21] = pc_init_val_o_21_sv2v_reg;
  assign pc_init_val_o[20] = pc_init_val_o_20_sv2v_reg;
  assign pc_init_val_o[19] = pc_init_val_o_19_sv2v_reg;
  assign pc_init_val_o[18] = pc_init_val_o_18_sv2v_reg;
  assign pc_init_val_o[17] = pc_init_val_o_17_sv2v_reg;
  assign pc_init_val_o[16] = pc_init_val_o_16_sv2v_reg;
  assign pc_init_val_o[15] = pc_init_val_o_15_sv2v_reg;
  assign pc_init_val_o[14] = pc_init_val_o_14_sv2v_reg;
  assign pc_init_val_o[13] = pc_init_val_o_13_sv2v_reg;
  assign pc_init_val_o[12] = pc_init_val_o_12_sv2v_reg;
  assign pc_init_val_o[11] = pc_init_val_o_11_sv2v_reg;
  assign pc_init_val_o[10] = pc_init_val_o_10_sv2v_reg;
  assign pc_init_val_o[9] = pc_init_val_o_9_sv2v_reg;
  assign pc_init_val_o[8] = pc_init_val_o_8_sv2v_reg;
  assign pc_init_val_o[7] = pc_init_val_o_7_sv2v_reg;
  assign pc_init_val_o[6] = pc_init_val_o_6_sv2v_reg;
  assign pc_init_val_o[5] = pc_init_val_o_5_sv2v_reg;
  assign pc_init_val_o[4] = pc_init_val_o_4_sv2v_reg;
  assign pc_init_val_o[3] = pc_init_val_o_3_sv2v_reg;
  assign pc_init_val_o[2] = pc_init_val_o_2_sv2v_reg;
  assign pc_init_val_o[1] = pc_init_val_o_1_sv2v_reg;
  assign pc_init_val_o[0] = pc_init_val_o_0_sv2v_reg;
  assign send_dmem_data_r = send_dmem_data_r_sv2v_reg;
  assign send_freeze_r = send_freeze_r_sv2v_reg;
  assign send_tgo_x_r = send_tgo_x_r_sv2v_reg;
  assign send_tgo_y_r = send_tgo_y_r_sv2v_reg;
  assign send_pc_init_val_r = send_pc_init_val_r_sv2v_reg;
  assign send_invalid_r = send_invalid_r_sv2v_reg;
  assign send_zero_r = send_zero_r_sv2v_reg;
  assign send_remote_interrupt_r = send_remote_interrupt_r_sv2v_reg;
  assign remote_dmem_addr_o[9] = addr_i[9];
  assign icache_pc_o[9] = remote_dmem_addr_o[9];
  assign remote_dmem_addr_o[8] = addr_i[8];
  assign icache_pc_o[8] = remote_dmem_addr_o[8];
  assign remote_dmem_addr_o[7] = addr_i[7];
  assign icache_pc_o[7] = remote_dmem_addr_o[7];
  assign remote_dmem_addr_o[6] = addr_i[6];
  assign icache_pc_o[6] = remote_dmem_addr_o[6];
  assign remote_dmem_addr_o[5] = addr_i[5];
  assign icache_pc_o[5] = remote_dmem_addr_o[5];
  assign remote_dmem_addr_o[4] = addr_i[4];
  assign icache_pc_o[4] = remote_dmem_addr_o[4];
  assign remote_dmem_addr_o[3] = addr_i[3];
  assign icache_pc_o[3] = remote_dmem_addr_o[3];
  assign remote_dmem_addr_o[2] = addr_i[2];
  assign icache_pc_o[2] = remote_dmem_addr_o[2];
  assign remote_dmem_addr_o[1] = addr_i[1];
  assign icache_pc_o[1] = remote_dmem_addr_o[1];
  assign remote_dmem_addr_o[0] = addr_i[0];
  assign icache_pc_o[0] = remote_dmem_addr_o[0];
  assign remote_dmem_mask_o[3] = mask_i[3];
  assign remote_dmem_mask_o[2] = mask_i[2];
  assign remote_dmem_mask_o[1] = mask_i[1];
  assign remote_dmem_mask_o[0] = mask_i[0];
  assign remote_dmem_data_o[31] = data_i[31];
  assign icache_instr_o[31] = remote_dmem_data_o[31];
  assign remote_dmem_data_o[30] = data_i[30];
  assign icache_instr_o[30] = remote_dmem_data_o[30];
  assign remote_dmem_data_o[29] = data_i[29];
  assign icache_instr_o[29] = remote_dmem_data_o[29];
  assign remote_dmem_data_o[28] = data_i[28];
  assign icache_instr_o[28] = remote_dmem_data_o[28];
  assign remote_dmem_data_o[27] = data_i[27];
  assign icache_instr_o[27] = remote_dmem_data_o[27];
  assign remote_dmem_data_o[26] = data_i[26];
  assign icache_instr_o[26] = remote_dmem_data_o[26];
  assign remote_dmem_data_o[25] = data_i[25];
  assign icache_instr_o[25] = remote_dmem_data_o[25];
  assign remote_dmem_data_o[24] = data_i[24];
  assign icache_instr_o[24] = remote_dmem_data_o[24];
  assign remote_dmem_data_o[23] = data_i[23];
  assign icache_instr_o[23] = remote_dmem_data_o[23];
  assign remote_dmem_data_o[22] = data_i[22];
  assign icache_instr_o[22] = remote_dmem_data_o[22];
  assign remote_dmem_data_o[21] = data_i[21];
  assign icache_instr_o[21] = remote_dmem_data_o[21];
  assign remote_dmem_data_o[20] = data_i[20];
  assign icache_instr_o[20] = remote_dmem_data_o[20];
  assign remote_dmem_data_o[19] = data_i[19];
  assign icache_instr_o[19] = remote_dmem_data_o[19];
  assign remote_dmem_data_o[18] = data_i[18];
  assign icache_instr_o[18] = remote_dmem_data_o[18];
  assign remote_dmem_data_o[17] = data_i[17];
  assign icache_instr_o[17] = remote_dmem_data_o[17];
  assign remote_dmem_data_o[16] = data_i[16];
  assign icache_instr_o[16] = remote_dmem_data_o[16];
  assign remote_dmem_data_o[15] = data_i[15];
  assign icache_instr_o[15] = remote_dmem_data_o[15];
  assign remote_dmem_data_o[14] = data_i[14];
  assign icache_instr_o[14] = remote_dmem_data_o[14];
  assign remote_dmem_data_o[13] = data_i[13];
  assign icache_instr_o[13] = remote_dmem_data_o[13];
  assign remote_dmem_data_o[12] = data_i[12];
  assign icache_instr_o[12] = remote_dmem_data_o[12];
  assign remote_dmem_data_o[11] = data_i[11];
  assign icache_instr_o[11] = remote_dmem_data_o[11];
  assign remote_dmem_data_o[10] = data_i[10];
  assign icache_instr_o[10] = remote_dmem_data_o[10];
  assign remote_dmem_data_o[9] = data_i[9];
  assign icache_instr_o[9] = remote_dmem_data_o[9];
  assign remote_dmem_data_o[8] = data_i[8];
  assign icache_instr_o[8] = remote_dmem_data_o[8];
  assign remote_dmem_data_o[7] = data_i[7];
  assign icache_instr_o[7] = remote_dmem_data_o[7];
  assign remote_dmem_data_o[6] = data_i[6];
  assign icache_instr_o[6] = remote_dmem_data_o[6];
  assign remote_dmem_data_o[5] = data_i[5];
  assign icache_instr_o[5] = remote_dmem_data_o[5];
  assign remote_dmem_data_o[4] = data_i[4];
  assign icache_instr_o[4] = remote_dmem_data_o[4];
  assign remote_dmem_data_o[3] = data_i[3];
  assign icache_instr_o[3] = remote_dmem_data_o[3];
  assign remote_dmem_data_o[2] = data_i[2];
  assign icache_instr_o[2] = remote_dmem_data_o[2];
  assign remote_dmem_data_o[1] = data_i[1];
  assign icache_instr_o[1] = remote_dmem_data_o[1];
  assign remote_dmem_data_o[0] = data_i[0];
  assign icache_instr_o[0] = remote_dmem_data_o[0];
  assign icache_pc_o_21_ = addr_i[21];
  assign icache_pc_o[21] = icache_pc_o_21_;
  assign icache_pc_o_20_ = addr_i[20];
  assign icache_pc_o[20] = icache_pc_o_20_;
  assign icache_pc_o_19_ = addr_i[19];
  assign icache_pc_o[19] = icache_pc_o_19_;
  assign icache_pc_o_18_ = addr_i[18];
  assign icache_pc_o[18] = icache_pc_o_18_;
  assign icache_pc_o_17_ = addr_i[17];
  assign icache_pc_o[17] = icache_pc_o_17_;
  assign icache_pc_o_16_ = addr_i[16];
  assign icache_pc_o[16] = icache_pc_o_16_;
  assign icache_pc_o_15_ = addr_i[15];
  assign icache_pc_o[15] = icache_pc_o_15_;
  assign icache_pc_o_14_ = addr_i[14];
  assign icache_pc_o[14] = icache_pc_o_14_;
  assign icache_pc_o_13_ = addr_i[13];
  assign icache_pc_o[13] = icache_pc_o_13_;
  assign icache_pc_o_12_ = addr_i[12];
  assign icache_pc_o[12] = icache_pc_o_12_;
  assign icache_pc_o_11_ = addr_i[11];
  assign icache_pc_o[11] = icache_pc_o_11_;
  assign icache_pc_o_10_ = addr_i[10];
  assign icache_pc_o[10] = icache_pc_o_10_;

  load_packer
  lp0
  (
    .mem_data_i(remote_dmem_data_i),
    .unsigned_load_i(load_info_r_is_unsigned_op_),
    .byte_load_i(load_info_r_is_byte_op_),
    .hex_load_i(load_info_r_is_hex_op_),
    .part_sel_i({ load_info_r_part_sel__1_, load_info_r_part_sel__0_ }),
    .load_data_o(load_data_lo)
  );

  assign N136 = reset_i | N7;
  assign N182 = ~icache_pc_o_13_;
  assign N183 = ~icache_pc_o_12_;
  assign N184 = ~icache_pc_o_11_;
  assign N185 = ~icache_pc_o_10_;
  assign N186 = ~remote_dmem_addr_o[9];
  assign N187 = ~remote_dmem_addr_o[8];
  assign N188 = ~remote_dmem_addr_o[7];
  assign N189 = ~remote_dmem_addr_o[6];
  assign N190 = ~remote_dmem_addr_o[5];
  assign N191 = ~remote_dmem_addr_o[4];
  assign N192 = ~remote_dmem_addr_o[3];
  assign N193 = ~remote_dmem_addr_o[2];
  assign N194 = ~remote_dmem_addr_o[1];
  assign N195 = ~remote_dmem_addr_o[0];
  assign N196 = icache_pc_o_21_ | N292;
  assign N197 = icache_pc_o_20_ | N196;
  assign N198 = icache_pc_o_19_ | N197;
  assign N199 = icache_pc_o_18_ | N198;
  assign N200 = icache_pc_o_17_ | N199;
  assign N201 = icache_pc_o_16_ | N200;
  assign N202 = icache_pc_o_15_ | N201;
  assign N203 = icache_pc_o_14_ | N202;
  assign N204 = N182 | N203;
  assign N205 = N183 | N204;
  assign N206 = N184 | N205;
  assign N207 = N185 | N206;
  assign N208 = N186 | N207;
  assign N209 = N187 | N208;
  assign N210 = N188 | N209;
  assign N211 = N189 | N210;
  assign N212 = N190 | N211;
  assign N213 = N191 | N212;
  assign N214 = N192 | N213;
  assign N215 = N193 | N214;
  assign N216 = N194 | N215;
  assign N217 = N195 | N216;
  assign N218 = ~N217;
  assign N219 = icache_pc_o_13_ | icache_pc_o_14_;
  assign N220 = icache_pc_o_12_ | N219;
  assign N221 = icache_pc_o_11_ | N220;
  assign N222 = icache_pc_o_10_ | N221;
  assign N223 = remote_dmem_addr_o[9] | N222;
  assign N224 = remote_dmem_addr_o[8] | N223;
  assign N225 = remote_dmem_addr_o[7] | N224;
  assign N226 = remote_dmem_addr_o[6] | N225;
  assign N227 = remote_dmem_addr_o[5] | N226;
  assign N228 = remote_dmem_addr_o[4] | N227;
  assign N229 = remote_dmem_addr_o[3] | N228;
  assign N230 = remote_dmem_addr_o[2] | N229;
  assign N231 = N194 | N230;
  assign N232 = N195 | N231;
  assign N233 = ~N232;
  assign N234 = icache_pc_o_13_ | icache_pc_o_14_;
  assign N235 = icache_pc_o_12_ | N234;
  assign N236 = icache_pc_o_11_ | N235;
  assign N237 = icache_pc_o_10_ | N236;
  assign N238 = remote_dmem_addr_o[9] | N237;
  assign N239 = remote_dmem_addr_o[8] | N238;
  assign N240 = remote_dmem_addr_o[7] | N239;
  assign N241 = remote_dmem_addr_o[6] | N240;
  assign N242 = remote_dmem_addr_o[5] | N241;
  assign N243 = remote_dmem_addr_o[4] | N242;
  assign N244 = remote_dmem_addr_o[3] | N243;
  assign N245 = remote_dmem_addr_o[2] | N244;
  assign N246 = N194 | N245;
  assign N247 = remote_dmem_addr_o[0] | N246;
  assign N248 = ~N247;
  assign N249 = icache_pc_o_13_ | icache_pc_o_14_;
  assign N250 = icache_pc_o_12_ | N249;
  assign N251 = icache_pc_o_11_ | N250;
  assign N252 = icache_pc_o_10_ | N251;
  assign N253 = remote_dmem_addr_o[9] | N252;
  assign N254 = remote_dmem_addr_o[8] | N253;
  assign N255 = remote_dmem_addr_o[7] | N254;
  assign N256 = remote_dmem_addr_o[6] | N255;
  assign N257 = remote_dmem_addr_o[5] | N256;
  assign N258 = remote_dmem_addr_o[4] | N257;
  assign N259 = remote_dmem_addr_o[3] | N258;
  assign N260 = remote_dmem_addr_o[2] | N259;
  assign N261 = remote_dmem_addr_o[1] | N260;
  assign N262 = N195 | N261;
  assign N263 = ~N262;
  assign N264 = icache_pc_o_13_ | icache_pc_o_14_;
  assign N265 = icache_pc_o_12_ | N264;
  assign N266 = icache_pc_o_11_ | N265;
  assign N267 = icache_pc_o_10_ | N266;
  assign N268 = remote_dmem_addr_o[9] | N267;
  assign N269 = remote_dmem_addr_o[8] | N268;
  assign N270 = remote_dmem_addr_o[7] | N269;
  assign N271 = remote_dmem_addr_o[6] | N270;
  assign N272 = remote_dmem_addr_o[5] | N271;
  assign N273 = remote_dmem_addr_o[4] | N272;
  assign N274 = remote_dmem_addr_o[3] | N273;
  assign N275 = remote_dmem_addr_o[2] | N274;
  assign N276 = remote_dmem_addr_o[1] | N275;
  assign N277 = remote_dmem_addr_o[0] | N276;
  assign N278 = ~N277;
  assign N279 = icache_pc_o_21_ | N292;
  assign N280 = icache_pc_o_20_ | N279;
  assign N281 = icache_pc_o_19_ | N280;
  assign N282 = icache_pc_o_18_ | N281;
  assign N283 = icache_pc_o_17_ | N282;
  assign N284 = icache_pc_o_16_ | N283;
  assign N285 = icache_pc_o_15_ | N284;
  assign N286 = icache_pc_o_14_ | N285;
  assign N287 = icache_pc_o_13_ | N286;
  assign N288 = icache_pc_o_12_ | N287;
  assign N289 = icache_pc_o_11_ | N288;
  assign N290 = icache_pc_o_10_ | N289;
  assign N291 = ~N290;
  assign N292 = addr_i[22] | N303;
  assign N293 = icache_pc_o_21_ | N292;
  assign N294 = icache_pc_o_20_ | N293;
  assign N295 = icache_pc_o_19_ | N294;
  assign N296 = icache_pc_o_18_ | N295;
  assign N297 = icache_pc_o_17_ | N296;
  assign N298 = icache_pc_o_16_ | N297;
  assign N299 = ~N298;
  assign N300 = addr_i[26] | addr_i[27];
  assign N301 = addr_i[25] | N300;
  assign N302 = addr_i[24] | N301;
  assign N303 = addr_i[23] | N302;
  assign N304 = ~N303;
  assign N23 = (N0)? 1'b1 : 
               (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N0 = N291;
  assign N1 = N290;
  assign N2 = 1'b0;
  assign N24 = (N0)? remote_dmem_yumi_i : 
               (N96)? icache_yumi_i : 
               (N99)? 1'b1 : 
               (N101)? 1'b1 : 
               (N103)? 1'b1 : 
               (N105)? 1'b1 : 
               (N107)? 1'b1 : 
               (N21)? 1'b1 : 1'b0;
  assign N25 = (N0)? remote_dmem_yumi_i : 
               (N96)? icache_yumi_i : 
               (N99)? 1'b1 : 
               (N101)? 1'b1 : 
               (N103)? 1'b1 : 
               (N105)? 1'b1 : 
               (N107)? 1'b1 : 
               (N21)? 1'b0 : 1'b0;
  assign N27 = (N0)? 1'b0 : 
               (N96)? 1'b1 : 
               (N26)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign { N33, N32, N31 } = (N103)? remote_dmem_data_o[2:0] : 
                             (N30)? tgo_y_o : 1'b0;
  assign { N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35 } = (N103)? pc_init_val_o : 
                                                                                                                            (N105)? remote_dmem_data_o[21:0] : 
                                                                                                                            (N34)? pc_init_val_o : 1'b0;
  assign N57 = (N0)? 1'b0 : 
               (N96)? 1'b0 : 
               (N99)? 1'b0 : 
               (N101)? 1'b0 : 
               (N103)? 1'b0 : 
               (N105)? 1'b0 : 
               (N107)? N22 : 
               (N21)? 1'b0 : 1'b0;
  assign N58 = (N0)? 1'b0 : 
               (N96)? 1'b0 : 
               (N99)? 1'b0 : 
               (N101)? 1'b0 : 
               (N103)? 1'b0 : 
               (N105)? 1'b0 : 
               (N107)? remote_dmem_data_o[0] : 
               (N21)? 1'b0 : 1'b0;
  assign N59 = (N0)? 1'b0 : 
               (N96)? 1'b0 : 
               (N99)? 1'b0 : 
               (N101)? 1'b0 : 
               (N103)? 1'b0 : 
               (N105)? 1'b0 : 
               (N107)? 1'b0 : 
               (N21)? 1'b1 : 1'b0;
  assign N61 = (N3)? N59 : 
               (N81)? 1'b0 : 
               (N83)? 1'b0 : 
               (N86)? 1'b0 : 
               (N89)? 1'b0 : 
               (N92)? 1'b0 : 
               (N95)? 1'b0 : 
               (N14)? 1'b1 : 1'b0;
  assign N3 = w_i;
  assign N63 = (N3)? N23 : 
               (N81)? 1'b1 : 
               (N62)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N65 = (N3)? N23 : 
               (N64)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N66 = (N3)? N24 : 
               (N81)? remote_dmem_yumi_i : 
               (N83)? 1'b1 : 
               (N86)? 1'b1 : 
               (N89)? 1'b1 : 
               (N92)? 1'b1 : 
               (N95)? 1'b1 : 
               (N14)? 1'b1 : 1'b0;
  assign N67 = (N3)? N25 : 
               (N64)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N68 = (N3)? N27 : 
               (N64)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N69 = (N3)? N57 : 
               (N64)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N70 = (N3)? N58 : 
               (N64)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N71 = (N3)? 1'b0 : 
               (N81)? remote_dmem_yumi_i : 
               (N62)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N73 = (N3)? 1'b0 : 
               (N81)? 1'b0 : 
               (N83)? 1'b1 : 
               (N72)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N75 = (N3)? 1'b0 : 
               (N81)? 1'b0 : 
               (N83)? 1'b0 : 
               (N86)? 1'b1 : 
               (N74)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N77 = (N3)? 1'b0 : 
               (N81)? 1'b0 : 
               (N83)? 1'b0 : 
               (N86)? 1'b0 : 
               (N89)? 1'b1 : 
               (N76)? 1'b0 : 
               (N2)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N79 = (N3)? 1'b0 : 
               (N81)? 1'b0 : 
               (N83)? 1'b0 : 
               (N86)? 1'b0 : 
               (N89)? 1'b0 : 
               (N92)? 1'b1 : 
               (N78)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N80 = (N3)? 1'b0 : 
               (N81)? 1'b0 : 
               (N83)? 1'b0 : 
               (N86)? 1'b0 : 
               (N89)? 1'b0 : 
               (N92)? 1'b0 : 
               (N95)? 1'b1 : 
               (N14)? 1'b0 : 1'b0;
  assign remote_dmem_v_o = (N4)? N63 : 
                           (N5)? 1'b0 : 1'b0;
  assign N4 = v_i;
  assign N5 = N7;
  assign remote_dmem_w_o = (N4)? N65 : 
                           (N5)? 1'b0 : 1'b0;
  assign yumi_o = (N4)? N66 : 
                  (N5)? 1'b0 : 1'b0;
  assign icache_v_o = (N4)? N68 : 
                      (N5)? 1'b0 : 1'b0;
  assign remote_interrupt_clear_o = (N4)? N69 : 
                                    (N5)? 1'b0 : 1'b0;
  assign remote_interrupt_set_o = (N4)? N70 : 
                                  (N5)? 1'b0 : 1'b0;
  assign returning_data_o = (N6)? load_data_lo : 
                            (N117)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, freeze_o } : 
                            (N120)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tgo_x_o } : 
                            (N123)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tgo_y_o } : 
                            (N126)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, pc_init_val_o } : 
                            (N129)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N132)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                            (N135)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, remote_interrupt_pending_bit_i } : 
                            (N115)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = send_dmem_data_r;
  assign is_icache_addr = addr_i[22] & N304;
  assign is_csr_addr = icache_pc_o_15_ & N299;
  assign is_freeze_addr = is_csr_addr & N278;
  assign is_tgo_x_addr = is_csr_addr & N263;
  assign is_tgo_y_addr = is_csr_addr & N248;
  assign is_pc_init_val_addr = is_csr_addr & N233;
  assign N7 = ~v_i;
  assign N8 = N291 | w_i;
  assign N9 = is_freeze_addr | N8;
  assign N10 = is_tgo_x_addr | N9;
  assign N11 = is_tgo_y_addr | N10;
  assign N12 = is_pc_init_val_addr | N11;
  assign N13 = N218 | N12;
  assign N14 = ~N13;
  assign N15 = is_icache_addr | N291;
  assign N16 = is_freeze_addr | N15;
  assign N17 = is_tgo_x_addr | N16;
  assign N18 = is_tgo_y_addr | N17;
  assign N19 = is_pc_init_val_addr | N18;
  assign N20 = N218 | N19;
  assign N21 = ~N20;
  assign N22 = ~remote_dmem_data_o[0];
  assign N26 = ~N15;
  assign N28 = ~N16;
  assign N29 = ~N17;
  assign N30 = ~N18;
  assign N34 = ~N19;
  assign N60 = ~remote_dmem_yumi_i;
  assign N62 = ~N8;
  assign N64 = ~w_i;
  assign N72 = ~N9;
  assign N74 = ~N10;
  assign N76 = ~N11;
  assign N78 = ~N12;
  assign N81 = N291 & N64;
  assign N82 = N64 & N290;
  assign N83 = is_freeze_addr & N82;
  assign N84 = ~is_freeze_addr;
  assign N85 = N82 & N84;
  assign N86 = is_tgo_x_addr & N85;
  assign N87 = ~is_tgo_x_addr;
  assign N88 = N85 & N87;
  assign N89 = is_tgo_y_addr & N88;
  assign N90 = ~is_tgo_y_addr;
  assign N91 = N88 & N90;
  assign N92 = is_pc_init_val_addr & N91;
  assign N93 = ~is_pc_init_val_addr;
  assign N94 = N91 & N93;
  assign N95 = N218 & N94;
  assign N96 = is_icache_addr & N290;
  assign N97 = ~is_icache_addr;
  assign N98 = N290 & N97;
  assign N99 = is_freeze_addr & N98;
  assign N100 = N98 & N84;
  assign N101 = is_tgo_x_addr & N100;
  assign N102 = N100 & N87;
  assign N103 = is_tgo_y_addr & N102;
  assign N104 = N102 & N90;
  assign N105 = is_pc_init_val_addr & N104;
  assign N106 = N104 & N93;
  assign N107 = N218 & N106;
  assign returning_data_v_o = N310 | send_remote_interrupt_r;
  assign N310 = N309 | send_zero_r;
  assign N309 = N308 | send_invalid_r;
  assign N308 = N307 | send_pc_init_val_r;
  assign N307 = N306 | send_tgo_y_r;
  assign N306 = N305 | send_tgo_x_r;
  assign N305 = send_dmem_data_r | send_freeze_r;
  assign N108 = send_freeze_r | send_dmem_data_r;
  assign N109 = send_tgo_x_r | N108;
  assign N110 = send_tgo_y_r | N109;
  assign N111 = send_pc_init_val_r | N110;
  assign N112 = send_zero_r | N111;
  assign N113 = send_invalid_r | N112;
  assign N114 = send_remote_interrupt_r | N113;
  assign N115 = ~N114;
  assign N116 = ~send_dmem_data_r;
  assign N117 = send_freeze_r & N116;
  assign N118 = ~send_freeze_r;
  assign N119 = N116 & N118;
  assign N120 = send_tgo_x_r & N119;
  assign N121 = ~send_tgo_x_r;
  assign N122 = N119 & N121;
  assign N123 = send_tgo_y_r & N122;
  assign N124 = ~send_tgo_y_r;
  assign N125 = N122 & N124;
  assign N126 = send_pc_init_val_r & N125;
  assign N127 = ~send_pc_init_val_r;
  assign N128 = N125 & N127;
  assign N129 = send_zero_r & N128;
  assign N130 = ~send_zero_r;
  assign N131 = N128 & N130;
  assign N132 = send_invalid_r & N131;
  assign N133 = ~send_invalid_r;
  assign N134 = N131 & N133;
  assign N135 = send_remote_interrupt_r & N134;
  assign N137 = w_i & v_i;
  assign N138 = N81 & v_i;
  assign N139 = N60 & N138;
  assign N140 = N137 | N139;
  assign N141 = N62 & v_i;
  assign N142 = N140 | N141;
  assign N143 = N142 | N7;
  assign N144 = ~N143;
  assign N145 = w_i & v_i;
  assign N146 = N145 | N139;
  assign N147 = N146 | N141;
  assign N148 = N147 | N7;
  assign N149 = ~N148;
  assign N150 = N291 & N145;
  assign N151 = N96 & N145;
  assign N152 = N150 | N151;
  assign N153 = N28 & N145;
  assign N154 = N152 | N153;
  assign N155 = N64 & v_i;
  assign N156 = N154 | N155;
  assign N157 = N156 | N7;
  assign N158 = ~N157;
  assign N159 = N99 & N145;
  assign N160 = N152 | N159;
  assign N161 = N29 & N145;
  assign N162 = N160 | N161;
  assign N163 = N162 | N155;
  assign N164 = N163 | N7;
  assign N165 = ~N164;
  assign N166 = N96 & N137;
  assign N167 = N150 | N166;
  assign N168 = N99 & N137;
  assign N169 = N167 | N168;
  assign N170 = N101 & N137;
  assign N171 = N169 | N170;
  assign N172 = N171 | N155;
  assign N173 = N172 | N7;
  assign N174 = ~N173;
  assign N175 = N291 & N137;
  assign N176 = N175 | N166;
  assign N177 = N176 | N168;
  assign N178 = N177 | N170;
  assign N179 = N178 | N155;
  assign N180 = N179 | N7;
  assign N181 = ~N180;

  always @(posedge clk_i) begin
    if(reset_i) begin
      load_info_r_is_unsigned_op__sv2v_reg <= 1'b0;
    end else if(N144) begin
      load_info_r_is_unsigned_op__sv2v_reg <= load_info_i[4];
    end 
    if(reset_i) begin
      load_info_r_is_byte_op__sv2v_reg <= 1'b0;
      load_info_r_is_hex_op__sv2v_reg <= 1'b0;
      load_info_r_part_sel__1__sv2v_reg <= 1'b0;
      load_info_r_part_sel__0__sv2v_reg <= 1'b0;
    end else if(N149) begin
      load_info_r_is_byte_op__sv2v_reg <= load_info_i[3];
      load_info_r_is_hex_op__sv2v_reg <= load_info_i[2];
      load_info_r_part_sel__1__sv2v_reg <= load_info_i[1];
      load_info_r_part_sel__0__sv2v_reg <= load_info_i[0];
    end 
    if(reset_i) begin
      freeze_o_sv2v_reg <= 1'b1;
    end else if(N158) begin
      freeze_o_sv2v_reg <= remote_dmem_data_o[0];
    end 
    if(reset_i) begin
      tgo_x_o_3_sv2v_reg <= 1'b0;
      tgo_x_o_2_sv2v_reg <= 1'b0;
      tgo_x_o_1_sv2v_reg <= 1'b0;
      tgo_x_o_0_sv2v_reg <= 1'b0;
    end else if(N165) begin
      tgo_x_o_3_sv2v_reg <= remote_dmem_data_o[3];
      tgo_x_o_2_sv2v_reg <= remote_dmem_data_o[2];
      tgo_x_o_1_sv2v_reg <= remote_dmem_data_o[1];
      tgo_x_o_0_sv2v_reg <= remote_dmem_data_o[0];
    end 
    if(reset_i) begin
      tgo_y_o_2_sv2v_reg <= 1'b0;
    end else if(N174) begin
      tgo_y_o_2_sv2v_reg <= N33;
    end 
    if(reset_i) begin
      tgo_y_o_1_sv2v_reg <= 1'b0;
      tgo_y_o_0_sv2v_reg <= 1'b0;
      pc_init_val_o_21_sv2v_reg <= 1'b0;
      pc_init_val_o_20_sv2v_reg <= 1'b0;
      pc_init_val_o_19_sv2v_reg <= 1'b0;
      pc_init_val_o_18_sv2v_reg <= 1'b0;
      pc_init_val_o_17_sv2v_reg <= 1'b0;
      pc_init_val_o_16_sv2v_reg <= 1'b0;
      pc_init_val_o_15_sv2v_reg <= 1'b0;
      pc_init_val_o_14_sv2v_reg <= 1'b0;
      pc_init_val_o_13_sv2v_reg <= 1'b0;
      pc_init_val_o_12_sv2v_reg <= 1'b0;
      pc_init_val_o_11_sv2v_reg <= 1'b0;
      pc_init_val_o_10_sv2v_reg <= 1'b0;
      pc_init_val_o_9_sv2v_reg <= 1'b0;
      pc_init_val_o_8_sv2v_reg <= 1'b0;
      pc_init_val_o_7_sv2v_reg <= 1'b0;
      pc_init_val_o_6_sv2v_reg <= 1'b0;
      pc_init_val_o_5_sv2v_reg <= 1'b0;
      pc_init_val_o_4_sv2v_reg <= 1'b0;
      pc_init_val_o_3_sv2v_reg <= 1'b0;
      pc_init_val_o_2_sv2v_reg <= 1'b0;
      pc_init_val_o_1_sv2v_reg <= 1'b0;
      pc_init_val_o_0_sv2v_reg <= 1'b0;
    end else if(N181) begin
      tgo_y_o_1_sv2v_reg <= N32;
      tgo_y_o_0_sv2v_reg <= N31;
      pc_init_val_o_21_sv2v_reg <= N56;
      pc_init_val_o_20_sv2v_reg <= N55;
      pc_init_val_o_19_sv2v_reg <= N54;
      pc_init_val_o_18_sv2v_reg <= N53;
      pc_init_val_o_17_sv2v_reg <= N52;
      pc_init_val_o_16_sv2v_reg <= N51;
      pc_init_val_o_15_sv2v_reg <= N50;
      pc_init_val_o_14_sv2v_reg <= N49;
      pc_init_val_o_13_sv2v_reg <= N48;
      pc_init_val_o_12_sv2v_reg <= N47;
      pc_init_val_o_11_sv2v_reg <= N46;
      pc_init_val_o_10_sv2v_reg <= N45;
      pc_init_val_o_9_sv2v_reg <= N44;
      pc_init_val_o_8_sv2v_reg <= N43;
      pc_init_val_o_7_sv2v_reg <= N42;
      pc_init_val_o_6_sv2v_reg <= N41;
      pc_init_val_o_5_sv2v_reg <= N40;
      pc_init_val_o_4_sv2v_reg <= N39;
      pc_init_val_o_3_sv2v_reg <= N38;
      pc_init_val_o_2_sv2v_reg <= N37;
      pc_init_val_o_1_sv2v_reg <= N36;
      pc_init_val_o_0_sv2v_reg <= N35;
    end 
    if(N136) begin
      send_dmem_data_r_sv2v_reg <= 1'b0;
      send_freeze_r_sv2v_reg <= 1'b0;
      send_tgo_x_r_sv2v_reg <= 1'b0;
      send_tgo_y_r_sv2v_reg <= 1'b0;
      send_pc_init_val_r_sv2v_reg <= 1'b0;
      send_invalid_r_sv2v_reg <= 1'b0;
      send_zero_r_sv2v_reg <= 1'b0;
      send_remote_interrupt_r_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      send_dmem_data_r_sv2v_reg <= N71;
      send_freeze_r_sv2v_reg <= N73;
      send_tgo_x_r_sv2v_reg <= N75;
      send_tgo_y_r_sv2v_reg <= N77;
      send_pc_init_val_r_sv2v_reg <= N79;
      send_invalid_r_sv2v_reg <= N61;
      send_zero_r_sv2v_reg <= N67;
      send_remote_interrupt_r_sv2v_reg <= N80;
    end 
  end


endmodule



module bsg_manycore_dram_hash_function_data_width_p32_addr_width_p28_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_x_subcord_width_p4_y_subcord_width_p3_num_vcache_rows_p1
(
  eva_i,
  pod_x_i,
  pod_y_i,
  epa_o,
  x_cord_o,
  y_cord_o
);

  input [31:0] eva_i;
  input [2:0] pod_x_i;
  input [3:0] pod_y_i;
  output [27:0] epa_o;
  output [6:0] x_cord_o;
  output [6:0] y_cord_o;
  wire [27:0] epa_o;
  wire [6:0] x_cord_o,y_cord_o;
  wire N0,epa_o_23_,epa_o_22_,epa_o_21_,epa_o_20_,epa_o_19_,epa_o_18_,epa_o_17_,
  epa_o_16_,epa_o_15_,epa_o_14_,epa_o_13_,epa_o_12_,epa_o_11_,epa_o_10_,epa_o_9_,
  epa_o_8_,epa_o_7_,epa_o_6_,epa_o_5_,epa_o_4_,epa_o_3_,epa_o_2_,epa_o_1_,epa_o_0_,N1,N2,
  N3,N4,N5,N6,N7,N8,N9;
  assign epa_o[24] = 1'b0;
  assign epa_o[25] = 1'b0;
  assign epa_o[26] = 1'b0;
  assign epa_o[27] = 1'b0;
  assign epa_o_23_ = eva_i[30];
  assign epa_o[23] = epa_o_23_;
  assign epa_o_22_ = eva_i[24];
  assign epa_o[22] = epa_o_22_;
  assign epa_o_21_ = eva_i[23];
  assign epa_o[21] = epa_o_21_;
  assign epa_o_20_ = eva_i[22];
  assign epa_o[20] = epa_o_20_;
  assign epa_o_19_ = eva_i[21];
  assign epa_o[19] = epa_o_19_;
  assign epa_o_18_ = eva_i[20];
  assign epa_o[18] = epa_o_18_;
  assign epa_o_17_ = eva_i[19];
  assign epa_o[17] = epa_o_17_;
  assign epa_o_16_ = eva_i[18];
  assign epa_o[16] = epa_o_16_;
  assign epa_o_15_ = eva_i[17];
  assign epa_o[15] = epa_o_15_;
  assign epa_o_14_ = eva_i[16];
  assign epa_o[14] = epa_o_14_;
  assign epa_o_13_ = eva_i[15];
  assign epa_o[13] = epa_o_13_;
  assign epa_o_12_ = eva_i[14];
  assign epa_o[12] = epa_o_12_;
  assign epa_o_11_ = eva_i[13];
  assign epa_o[11] = epa_o_11_;
  assign epa_o_10_ = eva_i[12];
  assign epa_o[10] = epa_o_10_;
  assign epa_o_9_ = eva_i[11];
  assign epa_o[9] = epa_o_9_;
  assign epa_o_8_ = eva_i[10];
  assign epa_o[8] = epa_o_8_;
  assign epa_o_7_ = eva_i[9];
  assign epa_o[7] = epa_o_7_;
  assign epa_o_6_ = eva_i[8];
  assign epa_o[6] = epa_o_6_;
  assign epa_o_5_ = eva_i[7];
  assign epa_o[5] = epa_o_5_;
  assign epa_o_4_ = eva_i[6];
  assign epa_o[4] = epa_o_4_;
  assign epa_o_3_ = eva_i[5];
  assign epa_o[3] = epa_o_3_;
  assign epa_o_2_ = eva_i[4];
  assign epa_o[2] = epa_o_2_;
  assign epa_o_1_ = eva_i[3];
  assign epa_o[1] = epa_o_1_;
  assign epa_o_0_ = eva_i[2];
  assign epa_o[0] = epa_o_0_;
  assign x_cord_o[6] = pod_x_i[2];
  assign x_cord_o[5] = pod_x_i[1];
  assign x_cord_o[4] = pod_x_i[0];
  assign x_cord_o[3] = eva_i[28];
  assign x_cord_o[2] = eva_i[27];
  assign x_cord_o[1] = eva_i[26];
  assign x_cord_o[0] = eva_i[25];
  assign { N5, N4, N3, N2 } = pod_y_i + 1'b1;
  assign { N9, N8, N7, N6 } = pod_y_i - 1'b1;
  assign y_cord_o[6:3] = (N0)? { N5, N4, N3, N2 } : 
                         (N1)? { N9, N8, N7, N6 } : 1'b0;
  assign N0 = eva_i[29];
  assign N1 = ~eva_i[29];
  assign y_cord_o[2] = ~eva_i[29];
  assign y_cord_o[1] = ~eva_i[29];
  assign y_cord_o[0] = ~eva_i[29];

endmodule



module bsg_manycore_eva_to_npa_data_width_p32_addr_width_p28_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_num_tiles_x_p16_num_tiles_y_p8_num_vcache_rows_p1_vcache_size_pinv_vcache_sets_pinv
(
  eva_i,
  tgo_x_i,
  tgo_y_i,
  pod_x_i,
  pod_y_i,
  x_cord_o,
  y_cord_o,
  epa_o,
  is_invalid_addr_o
);

  input [31:0] eva_i;
  input [3:0] tgo_x_i;
  input [2:0] tgo_y_i;
  input [2:0] pod_x_i;
  input [3:0] pod_y_i;
  output [6:0] x_cord_o;
  output [6:0] y_cord_o;
  output [27:0] epa_o;
  output is_invalid_addr_o;
  wire [6:0] x_cord_o,y_cord_o,dram_x_cord_lo,dram_y_cord_lo;
  wire [27:0] epa_o,dram_epa_lo;
  wire is_invalid_addr_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,N21,N22,N23;

  bsg_manycore_dram_hash_function_data_width_p32_addr_width_p28_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_x_subcord_width_p4_y_subcord_width_p3_num_vcache_rows_p1
  dram_hash
  (
    .eva_i(eva_i),
    .pod_x_i(pod_x_i),
    .pod_y_i(pod_y_i),
    .epa_o(dram_epa_lo),
    .x_cord_o(dram_x_cord_lo),
    .y_cord_o(dram_y_cord_lo)
  );

  assign N17 = ~eva_i[29];
  assign N18 = eva_i[30] | eva_i[31];
  assign N19 = N17 | N18;
  assign N20 = ~N19;
  assign N21 = ~eva_i[30];
  assign N22 = N21 | eva_i[31];
  assign N23 = ~N22;
  assign { N12, N11, N10, N9 } = eva_i[21:18] + tgo_x_i;
  assign { N8, N7, N6 } = eva_i[26:24] + tgo_y_i;
  assign y_cord_o = (N0)? dram_y_cord_lo : 
                    (N14)? eva_i[29:23] : 
                    (N16)? { pod_y_i, N8, N7, N6 } : 
                    (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N1;
  assign x_cord_o = (N0)? dram_x_cord_lo : 
                    (N14)? eva_i[22:16] : 
                    (N16)? { pod_x_i, N12, N11, N10, N9 } : 
                    (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign epa_o = (N0)? dram_epa_lo : 
                 (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, eva_i[15:2] } : 
                 (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, eva_i[17:2] } : 
                 (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign is_invalid_addr_o = (N0)? 1'b0 : 
                             (N14)? 1'b0 : 
                             (N16)? 1'b0 : 
                             (N4)? 1'b1 : 1'b0;
  assign N1 = eva_i[31];
  assign N2 = N23 | N1;
  assign N3 = N20 | N2;
  assign N4 = ~N3;
  assign N5 = N16;
  assign N13 = ~N1;
  assign N14 = N23 & N13;
  assign N15 = N13 & N22;
  assign N16 = N20 & N15;

endmodule



module network_tx_data_width_p32_addr_width_p28_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_num_vcache_rows_p1_vcache_size_pinv_vcache_sets_pinv_num_tiles_x_p16_num_tiles_y_p8_icache_entries_p1024_icache_tag_width_p12
(
  clk_i,
  reset_i,
  out_packet_o,
  out_v_o,
  out_credit_or_ready_i,
  returned_v_i,
  returned_data_i,
  returned_reg_id_i,
  returned_pkt_type_i,
  returned_fifo_full_i,
  returned_yumi_o,
  tgo_x_i,
  tgo_y_i,
  my_x_i,
  my_y_i,
  pod_x_i,
  pod_y_i,
  cfg_pod_x_i,
  cfg_pod_y_i,
  remote_req_i,
  remote_req_v_i,
  remote_req_credit_o,
  ifetch_v_o,
  ifetch_instr_o,
  float_remote_load_resp_rd_o,
  float_remote_load_resp_data_o,
  float_remote_load_resp_v_o,
  float_remote_load_resp_force_o,
  float_remote_load_resp_yumi_i,
  int_remote_load_resp_rd_o,
  int_remote_load_resp_data_o,
  int_remote_load_resp_v_o,
  int_remote_load_resp_force_o,
  int_remote_load_resp_yumi_i,
  invalid_eva_access_o
);

  output [96:0] out_packet_o;
  input [31:0] returned_data_i;
  input [4:0] returned_reg_id_i;
  input [1:0] returned_pkt_type_i;
  input [3:0] tgo_x_i;
  input [2:0] tgo_y_i;
  input [3:0] my_x_i;
  input [2:0] my_y_i;
  input [2:0] pod_x_i;
  input [3:0] pod_y_i;
  input [2:0] cfg_pod_x_i;
  input [3:0] cfg_pod_y_i;
  input [83:0] remote_req_i;
  output [31:0] ifetch_instr_o;
  output [4:0] float_remote_load_resp_rd_o;
  output [31:0] float_remote_load_resp_data_o;
  output [4:0] int_remote_load_resp_rd_o;
  output [31:0] int_remote_load_resp_data_o;
  input clk_i;
  input reset_i;
  input out_credit_or_ready_i;
  input returned_v_i;
  input returned_fifo_full_i;
  input remote_req_v_i;
  input float_remote_load_resp_yumi_i;
  input int_remote_load_resp_yumi_i;
  output out_v_o;
  output returned_yumi_o;
  output remote_req_credit_o;
  output ifetch_v_o;
  output float_remote_load_resp_v_o;
  output float_remote_load_resp_force_o;
  output int_remote_load_resp_v_o;
  output int_remote_load_resp_force_o;
  output invalid_eva_access_o;
  wire [96:0] out_packet_o;
  wire [31:0] ifetch_instr_o,float_remote_load_resp_data_o,int_remote_load_resp_data_o;
  wire [4:0] float_remote_load_resp_rd_o,int_remote_load_resp_rd_o;
  wire out_v_o,returned_yumi_o,remote_req_credit_o,ifetch_v_o,
  float_remote_load_resp_v_o,float_remote_load_resp_force_o,int_remote_load_resp_v_o,
  int_remote_load_resp_force_o,invalid_eva_access_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,out_packet_o_27_,
  out_packet_o_26_,out_packet_o_25_,out_packet_o_24_,out_packet_o_23_,
  out_packet_o_22_,out_packet_o_21_,out_packet_o_20_,out_packet_o_19_,out_packet_o_18_,
  out_packet_o_17_,out_packet_o_16_,out_packet_o_15_,out_packet_o_14_,is_invalid_addr_lo,
  _1_net__2_,_1_net__1_,_1_net__0_,_2_net__3_,_2_net__2_,_2_net__1_,_2_net__0_,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36;
  assign out_packet_o[66] = 1'b0;
  assign out_packet_o_27_ = pod_y_i[3];
  assign out_packet_o[27] = out_packet_o_27_;
  assign out_packet_o_26_ = pod_y_i[2];
  assign out_packet_o[26] = out_packet_o_26_;
  assign out_packet_o_25_ = pod_y_i[1];
  assign out_packet_o[25] = out_packet_o_25_;
  assign out_packet_o_24_ = pod_y_i[0];
  assign out_packet_o[24] = out_packet_o_24_;
  assign out_packet_o_23_ = my_y_i[2];
  assign out_packet_o[23] = out_packet_o_23_;
  assign out_packet_o_22_ = my_y_i[1];
  assign out_packet_o[22] = out_packet_o_22_;
  assign out_packet_o_21_ = my_y_i[0];
  assign out_packet_o[21] = out_packet_o_21_;
  assign out_packet_o_20_ = pod_x_i[2];
  assign out_packet_o[20] = out_packet_o_20_;
  assign out_packet_o_19_ = pod_x_i[1];
  assign out_packet_o[19] = out_packet_o_19_;
  assign out_packet_o_18_ = pod_x_i[0];
  assign out_packet_o[18] = out_packet_o_18_;
  assign out_packet_o_17_ = my_x_i[3];
  assign out_packet_o[17] = out_packet_o_17_;
  assign out_packet_o_16_ = my_x_i[2];
  assign out_packet_o[16] = out_packet_o_16_;
  assign out_packet_o_15_ = my_x_i[1];
  assign out_packet_o[15] = out_packet_o_15_;
  assign out_packet_o_14_ = my_x_i[0];
  assign out_packet_o[14] = out_packet_o_14_;
  assign remote_req_credit_o = out_credit_or_ready_i;
  assign ifetch_instr_o[31] = returned_data_i[31];
  assign float_remote_load_resp_data_o[31] = ifetch_instr_o[31];
  assign int_remote_load_resp_data_o[31] = ifetch_instr_o[31];
  assign ifetch_instr_o[30] = returned_data_i[30];
  assign float_remote_load_resp_data_o[30] = ifetch_instr_o[30];
  assign int_remote_load_resp_data_o[30] = ifetch_instr_o[30];
  assign ifetch_instr_o[29] = returned_data_i[29];
  assign float_remote_load_resp_data_o[29] = ifetch_instr_o[29];
  assign int_remote_load_resp_data_o[29] = ifetch_instr_o[29];
  assign ifetch_instr_o[28] = returned_data_i[28];
  assign float_remote_load_resp_data_o[28] = ifetch_instr_o[28];
  assign int_remote_load_resp_data_o[28] = ifetch_instr_o[28];
  assign ifetch_instr_o[27] = returned_data_i[27];
  assign float_remote_load_resp_data_o[27] = ifetch_instr_o[27];
  assign int_remote_load_resp_data_o[27] = ifetch_instr_o[27];
  assign ifetch_instr_o[26] = returned_data_i[26];
  assign float_remote_load_resp_data_o[26] = ifetch_instr_o[26];
  assign int_remote_load_resp_data_o[26] = ifetch_instr_o[26];
  assign ifetch_instr_o[25] = returned_data_i[25];
  assign float_remote_load_resp_data_o[25] = ifetch_instr_o[25];
  assign int_remote_load_resp_data_o[25] = ifetch_instr_o[25];
  assign ifetch_instr_o[24] = returned_data_i[24];
  assign float_remote_load_resp_data_o[24] = ifetch_instr_o[24];
  assign int_remote_load_resp_data_o[24] = ifetch_instr_o[24];
  assign ifetch_instr_o[23] = returned_data_i[23];
  assign float_remote_load_resp_data_o[23] = ifetch_instr_o[23];
  assign int_remote_load_resp_data_o[23] = ifetch_instr_o[23];
  assign ifetch_instr_o[22] = returned_data_i[22];
  assign float_remote_load_resp_data_o[22] = ifetch_instr_o[22];
  assign int_remote_load_resp_data_o[22] = ifetch_instr_o[22];
  assign ifetch_instr_o[21] = returned_data_i[21];
  assign float_remote_load_resp_data_o[21] = ifetch_instr_o[21];
  assign int_remote_load_resp_data_o[21] = ifetch_instr_o[21];
  assign ifetch_instr_o[20] = returned_data_i[20];
  assign float_remote_load_resp_data_o[20] = ifetch_instr_o[20];
  assign int_remote_load_resp_data_o[20] = ifetch_instr_o[20];
  assign ifetch_instr_o[19] = returned_data_i[19];
  assign float_remote_load_resp_data_o[19] = ifetch_instr_o[19];
  assign int_remote_load_resp_data_o[19] = ifetch_instr_o[19];
  assign ifetch_instr_o[18] = returned_data_i[18];
  assign float_remote_load_resp_data_o[18] = ifetch_instr_o[18];
  assign int_remote_load_resp_data_o[18] = ifetch_instr_o[18];
  assign ifetch_instr_o[17] = returned_data_i[17];
  assign float_remote_load_resp_data_o[17] = ifetch_instr_o[17];
  assign int_remote_load_resp_data_o[17] = ifetch_instr_o[17];
  assign ifetch_instr_o[16] = returned_data_i[16];
  assign float_remote_load_resp_data_o[16] = ifetch_instr_o[16];
  assign int_remote_load_resp_data_o[16] = ifetch_instr_o[16];
  assign ifetch_instr_o[15] = returned_data_i[15];
  assign float_remote_load_resp_data_o[15] = ifetch_instr_o[15];
  assign int_remote_load_resp_data_o[15] = ifetch_instr_o[15];
  assign ifetch_instr_o[14] = returned_data_i[14];
  assign float_remote_load_resp_data_o[14] = ifetch_instr_o[14];
  assign int_remote_load_resp_data_o[14] = ifetch_instr_o[14];
  assign ifetch_instr_o[13] = returned_data_i[13];
  assign float_remote_load_resp_data_o[13] = ifetch_instr_o[13];
  assign int_remote_load_resp_data_o[13] = ifetch_instr_o[13];
  assign ifetch_instr_o[12] = returned_data_i[12];
  assign float_remote_load_resp_data_o[12] = ifetch_instr_o[12];
  assign int_remote_load_resp_data_o[12] = ifetch_instr_o[12];
  assign ifetch_instr_o[11] = returned_data_i[11];
  assign float_remote_load_resp_data_o[11] = ifetch_instr_o[11];
  assign int_remote_load_resp_data_o[11] = ifetch_instr_o[11];
  assign ifetch_instr_o[10] = returned_data_i[10];
  assign float_remote_load_resp_data_o[10] = ifetch_instr_o[10];
  assign int_remote_load_resp_data_o[10] = ifetch_instr_o[10];
  assign ifetch_instr_o[9] = returned_data_i[9];
  assign float_remote_load_resp_data_o[9] = ifetch_instr_o[9];
  assign int_remote_load_resp_data_o[9] = ifetch_instr_o[9];
  assign ifetch_instr_o[8] = returned_data_i[8];
  assign float_remote_load_resp_data_o[8] = ifetch_instr_o[8];
  assign int_remote_load_resp_data_o[8] = ifetch_instr_o[8];
  assign ifetch_instr_o[7] = returned_data_i[7];
  assign float_remote_load_resp_data_o[7] = ifetch_instr_o[7];
  assign int_remote_load_resp_data_o[7] = ifetch_instr_o[7];
  assign ifetch_instr_o[6] = returned_data_i[6];
  assign float_remote_load_resp_data_o[6] = ifetch_instr_o[6];
  assign int_remote_load_resp_data_o[6] = ifetch_instr_o[6];
  assign ifetch_instr_o[5] = returned_data_i[5];
  assign float_remote_load_resp_data_o[5] = ifetch_instr_o[5];
  assign int_remote_load_resp_data_o[5] = ifetch_instr_o[5];
  assign ifetch_instr_o[4] = returned_data_i[4];
  assign float_remote_load_resp_data_o[4] = ifetch_instr_o[4];
  assign int_remote_load_resp_data_o[4] = ifetch_instr_o[4];
  assign ifetch_instr_o[3] = returned_data_i[3];
  assign float_remote_load_resp_data_o[3] = ifetch_instr_o[3];
  assign int_remote_load_resp_data_o[3] = ifetch_instr_o[3];
  assign ifetch_instr_o[2] = returned_data_i[2];
  assign float_remote_load_resp_data_o[2] = ifetch_instr_o[2];
  assign int_remote_load_resp_data_o[2] = ifetch_instr_o[2];
  assign ifetch_instr_o[1] = returned_data_i[1];
  assign float_remote_load_resp_data_o[1] = ifetch_instr_o[1];
  assign int_remote_load_resp_data_o[1] = ifetch_instr_o[1];
  assign ifetch_instr_o[0] = returned_data_i[0];
  assign float_remote_load_resp_data_o[0] = ifetch_instr_o[0];
  assign int_remote_load_resp_data_o[0] = ifetch_instr_o[0];
  assign int_remote_load_resp_rd_o[4] = returned_reg_id_i[4];
  assign float_remote_load_resp_rd_o[4] = int_remote_load_resp_rd_o[4];
  assign int_remote_load_resp_rd_o[3] = returned_reg_id_i[3];
  assign float_remote_load_resp_rd_o[3] = int_remote_load_resp_rd_o[3];
  assign int_remote_load_resp_rd_o[2] = returned_reg_id_i[2];
  assign float_remote_load_resp_rd_o[2] = int_remote_load_resp_rd_o[2];
  assign int_remote_load_resp_rd_o[1] = returned_reg_id_i[1];
  assign float_remote_load_resp_rd_o[1] = int_remote_load_resp_rd_o[1];
  assign int_remote_load_resp_rd_o[0] = returned_reg_id_i[0];
  assign float_remote_load_resp_rd_o[0] = int_remote_load_resp_rd_o[0];

  bsg_manycore_eva_to_npa_data_width_p32_addr_width_p28_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_num_tiles_x_p16_num_tiles_y_p8_num_vcache_rows_p1_vcache_size_pinv_vcache_sets_pinv
  eva2npa
  (
    .eva_i(remote_req_i[31:0]),
    .tgo_x_i(tgo_x_i),
    .tgo_y_i(tgo_y_i),
    .pod_x_i({ _1_net__2_, _1_net__1_, _1_net__0_ }),
    .pod_y_i({ _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ }),
    .x_cord_o(out_packet_o[6:0]),
    .y_cord_o(out_packet_o[13:7]),
    .epa_o(out_packet_o[96:69]),
    .is_invalid_addr_o(is_invalid_addr_lo)
  );

  assign N19 = N17 & N18;
  assign N20 = remote_req_i[81] | N18;
  assign N22 = N17 | remote_req_i[80];
  assign N24 = remote_req_i[81] & remote_req_i[80];
  assign N32 = returned_pkt_type_i[0] & returned_pkt_type_i[1];
  assign N33 = ~returned_pkt_type_i[1];
  assign N34 = returned_pkt_type_i[0] | N33;
  assign N35 = ~N34;
  assign { _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ } = (N0)? { out_packet_o_27_, out_packet_o_26_, out_packet_o_25_, out_packet_o_24_ } : 
                                                              (N11)? cfg_pod_y_i : 1'b0;
  assign N0 = remote_req_i[74];
  assign { _1_net__2_, _1_net__1_, _1_net__0_ } = (N0)? { out_packet_o_20_, out_packet_o_19_, out_packet_o_18_ } : 
                                                  (N11)? cfg_pod_x_i : 1'b0;
  assign out_packet_o[59:28] = (N1)? remote_req_i[63:32] : 
                               (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, remote_req_i[75:69] } : 1'b0;
  assign N1 = N12;
  assign out_packet_o[64:60] = (N2)? { 1'b0, remote_req_i[79:76] } : 
                               (N14)? remote_req_i[68:64] : 1'b0;
  assign N2 = remote_req_i[83];
  assign { N27, N26, N25 } = (N3)? { 1'b0, 1'b1, 1'b0 } : 
                             (N4)? { 1'b1, 1'b0, 1'b0 } : 
                             (N5)? { 1'b0, 1'b1, 1'b1 } : 
                             (N6)? { 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign N3 = N19;
  assign N4 = N21;
  assign N5 = N23;
  assign N6 = N24;
  assign { out_packet_o[68:67], out_packet_o[65:65] } = (N7)? { N27, N26, N25 } : 
                                                        (N29)? { 1'b0, 1'b0, 1'b1 } : 
                                                        (N16)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = remote_req_i[82];
  assign ifetch_v_o = (N8)? returned_v_i : 
                      (N9)? 1'b0 : 
                      (N10)? 1'b0 : 1'b0;
  assign N8 = N32;
  assign N9 = N35;
  assign N10 = N33;
  assign returned_yumi_o = (N8)? returned_v_i : 
                           (N9)? N30 : 
                           (N10)? N31 : 1'b0;
  assign float_remote_load_resp_v_o = (N8)? 1'b0 : 
                                      (N9)? returned_v_i : 
                                      (N10)? 1'b0 : 1'b0;
  assign float_remote_load_resp_force_o = (N8)? 1'b0 : 
                                          (N9)? returned_fifo_full_i : 
                                          (N10)? 1'b0 : 1'b0;
  assign int_remote_load_resp_v_o = (N8)? 1'b0 : 
                                    (N9)? 1'b0 : 
                                    (N10)? returned_v_i : 1'b0;
  assign int_remote_load_resp_force_o = (N8)? 1'b0 : 
                                        (N9)? 1'b0 : 
                                        (N10)? returned_fifo_full_i : 1'b0;
  assign N11 = ~remote_req_i[74];
  assign N12 = remote_req_i[83] | remote_req_i[82];
  assign N13 = ~N12;
  assign N14 = ~remote_req_i[83];
  assign N15 = remote_req_i[83] | remote_req_i[82];
  assign N16 = ~N15;
  assign N17 = ~remote_req_i[81];
  assign N18 = ~remote_req_i[80];
  assign N21 = ~N20;
  assign N23 = ~N22;
  assign N28 = ~remote_req_i[82];
  assign N29 = remote_req_i[83] & N28;
  assign out_v_o = remote_req_v_i & N36;
  assign N36 = ~is_invalid_addr_lo;
  assign invalid_eva_access_o = remote_req_v_i & is_invalid_addr_lo;
  assign N30 = float_remote_load_resp_yumi_i | returned_fifo_full_i;
  assign N31 = int_remote_load_resp_yumi_i | returned_fifo_full_i;

endmodule



module bsg_mem_1rw_sync_width_p46_els_p1024_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [45:0] data_i;
  input [9:0] addr_i;
  output [45:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [45:0] data_o;

//   fakeram130_1024x46 fakeram2
//	(
//	   data_o,
//  	 addr_i,
// 	  w_i,
// 	  data_i,
//  	 w_mask_in,
//  	 clk_i,
//  	 v_i
//	);

  hard_mem_1rw_d1024_w46_wrapper
  \macro.mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(w_i),
    .data_o(data_o)
   );


endmodule



module icache_icache_tag_width_p12_icache_entries_p1024
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  flush_i,
  w_pc_i,
  w_instr_i,
  pc_i,
  jalr_prediction_i,
  instr_o,
  pred_or_jump_addr_o,
  pc_r_o,
  icache_miss_o,
  icache_flush_r_o
);

  input [21:0] w_pc_i;
  input [31:0] w_instr_i;
  input [21:0] pc_i;
  input [21:0] jalr_prediction_i;
  output [31:0] instr_o;
  output [21:0] pred_or_jump_addr_o;
  output [21:0] pc_r_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  input flush_i;
  output icache_miss_o;
  output icache_flush_r_o;
  wire [31:0] instr_o;
  wire [21:0] pred_or_jump_addr_o,pc_r_o;
  wire icache_miss_o,icache_flush_r_o,N0,N1,N2,N3,N4,N5,icache_data_li_lower_cout_,
  icache_data_lo_lower_cout_,icache_data_lo_lower_sign_,icache_data_lo_tag__11_,
  icache_data_lo_tag__10_,icache_data_lo_tag__9_,icache_data_lo_tag__8_,
  icache_data_lo_tag__7_,icache_data_lo_tag__6_,icache_data_lo_tag__5_,icache_data_lo_tag__4_,
  icache_data_lo_tag__3_,icache_data_lo_tag__2_,icache_data_lo_tag__1_,
  icache_data_lo_tag__0_,N6,N7,write_branch_instr,write_jal_instr,branch_pc_lower_cout,
  jal_pc_lower_cout,N8,N9,injected_instr_0,N10,N11,N12,N13,N14,N15,sel_pc,sel_pc_p1,N16,N17,
  N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,
  N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,
  N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,
  N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  sv2v_dc_1,sv2v_dc_2;
  wire [9:0] icache_addr_li;
  wire [12:1] branch_pc_lower_res;
  wire [20:1] jal_pc_lower_res;
  wire [31:7] injected_instr;
  wire [10:0] branch_pc_high_out;
  wire [2:0] jal_pc_high_out;
  reg icache_flush_r_o_sv2v_reg,pc_r_o_21_sv2v_reg,pc_r_o_20_sv2v_reg,
  pc_r_o_19_sv2v_reg,pc_r_o_18_sv2v_reg,pc_r_o_17_sv2v_reg,pc_r_o_16_sv2v_reg,pc_r_o_15_sv2v_reg,
  pc_r_o_14_sv2v_reg,pc_r_o_13_sv2v_reg,pc_r_o_12_sv2v_reg,pc_r_o_11_sv2v_reg,
  pc_r_o_10_sv2v_reg,pc_r_o_9_sv2v_reg,pc_r_o_8_sv2v_reg,pc_r_o_7_sv2v_reg,
  pc_r_o_6_sv2v_reg,pc_r_o_5_sv2v_reg,pc_r_o_4_sv2v_reg,pc_r_o_3_sv2v_reg,pc_r_o_2_sv2v_reg,
  pc_r_o_1_sv2v_reg,pc_r_o_0_sv2v_reg;
  assign icache_flush_r_o = icache_flush_r_o_sv2v_reg;
  assign pc_r_o[21] = pc_r_o_21_sv2v_reg;
  assign pc_r_o[20] = pc_r_o_20_sv2v_reg;
  assign pc_r_o[19] = pc_r_o_19_sv2v_reg;
  assign pc_r_o[18] = pc_r_o_18_sv2v_reg;
  assign pc_r_o[17] = pc_r_o_17_sv2v_reg;
  assign pc_r_o[16] = pc_r_o_16_sv2v_reg;
  assign pc_r_o[15] = pc_r_o_15_sv2v_reg;
  assign pc_r_o[14] = pc_r_o_14_sv2v_reg;
  assign pc_r_o[13] = pc_r_o_13_sv2v_reg;
  assign pc_r_o[12] = pc_r_o_12_sv2v_reg;
  assign pc_r_o[11] = pc_r_o_11_sv2v_reg;
  assign pc_r_o[10] = pc_r_o_10_sv2v_reg;
  assign pc_r_o[9] = pc_r_o_9_sv2v_reg;
  assign pc_r_o[8] = pc_r_o_8_sv2v_reg;
  assign pc_r_o[7] = pc_r_o_7_sv2v_reg;
  assign pc_r_o[6] = pc_r_o_6_sv2v_reg;
  assign pc_r_o[5] = pc_r_o_5_sv2v_reg;
  assign pc_r_o[4] = pc_r_o_4_sv2v_reg;
  assign pc_r_o[3] = pc_r_o_3_sv2v_reg;
  assign pc_r_o[2] = pc_r_o_2_sv2v_reg;
  assign pc_r_o[1] = pc_r_o_1_sv2v_reg;
  assign pc_r_o[0] = pc_r_o_0_sv2v_reg;

  bsg_mem_1rw_sync_width_p46_els_p1024_latch_last_read_p1
  imem_0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ icache_data_li_lower_cout_, w_instr_i[31:31], w_pc_i[21:10], injected_instr, w_instr_i[6:1], injected_instr_0 }),
    .addr_i(icache_addr_li),
    .v_i(v_i),
    .w_i(w_i),
    .data_o({ icache_data_lo_lower_cout_, icache_data_lo_lower_sign_, icache_data_lo_tag__11_, icache_data_lo_tag__10_, icache_data_lo_tag__9_, icache_data_lo_tag__8_, icache_data_lo_tag__7_, icache_data_lo_tag__6_, icache_data_lo_tag__5_, icache_data_lo_tag__4_, icache_data_lo_tag__3_, icache_data_lo_tag__2_, icache_data_lo_tag__1_, icache_data_lo_tag__0_, instr_o })
  );

  assign icache_miss_o = { icache_data_lo_tag__11_, icache_data_lo_tag__10_, icache_data_lo_tag__9_, icache_data_lo_tag__8_, icache_data_lo_tag__7_, icache_data_lo_tag__6_, icache_data_lo_tag__5_, icache_data_lo_tag__4_, icache_data_lo_tag__3_, icache_data_lo_tag__2_, icache_data_lo_tag__1_, icache_data_lo_tag__0_ } != pc_r_o[21:10];
  assign N52 = reset_i | N13;
  assign N53 = ~instr_o[6];
  assign N54 = ~instr_o[5];
  assign N55 = ~instr_o[2];
  assign N56 = ~instr_o[1];
  assign N57 = ~instr_o[0];
  assign N58 = N54 | N53;
  assign N59 = instr_o[4] | N58;
  assign N60 = instr_o[3] | N59;
  assign N61 = N55 | N60;
  assign N62 = N56 | N61;
  assign N63 = N57 | N62;
  assign N64 = ~N63;
  assign N65 = ~instr_o[3];
  assign N66 = N54 | N53;
  assign N67 = instr_o[4] | N66;
  assign N68 = N65 | N67;
  assign N69 = N55 | N68;
  assign N70 = N56 | N69;
  assign N71 = N57 | N70;
  assign N72 = ~N71;
  assign { branch_pc_lower_cout, branch_pc_lower_res, sv2v_dc_1 } = { w_instr_i[31:31], w_instr_i[7:7], w_instr_i[30:25], w_instr_i[11:8], 1'b0 } + { w_pc_i[10:0], 1'b0, 1'b0 };
  assign { jal_pc_lower_cout, jal_pc_lower_res, sv2v_dc_2 } = { w_instr_i[31:31], w_instr_i[19:12], w_instr_i[20:20], w_instr_i[30:21], 1'b0 } + { w_pc_i[18:0], 1'b0, 1'b0 };
  assign { N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33 } = pc_r_o[21:11] - 1'b1;
  assign { N46, N45, N44 } = pc_r_o[21:19] - 1'b1;
  assign { N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19 } = pc_r_o[21:11] + 1'b1;
  assign { N32, N31, N30 } = pc_r_o[21:19] + 1'b1;
  assign icache_addr_li = (N0)? w_pc_i[9:0] : 
                          (N7)? pc_i[9:0] : 1'b0;
  assign N0 = N6;
  assign { injected_instr, injected_instr_0 } = (N1)? { branch_pc_lower_res[12:12], branch_pc_lower_res[10:5], w_instr_i[24:12], branch_pc_lower_res[4:1], branch_pc_lower_res[11:11], w_instr_i[31:31] } : 
                                                (N11)? { jal_pc_lower_res[20:20], jal_pc_lower_res[10:1], jal_pc_lower_res[11:11], jal_pc_lower_res[19:12], w_instr_i[11:7], w_instr_i[0:0] } : 
                                                (N9)? { w_instr_i[31:7], w_instr_i[0:0] } : 1'b0;
  assign N1 = write_branch_instr;
  assign icache_data_li_lower_cout_ = (N1)? branch_pc_lower_cout : 
                                      (N2)? jal_pc_lower_cout : 1'b0;
  assign N2 = N12;
  assign N15 = (N3)? 1'b1 : 
               (N14)? 1'b0 : 1'b0;
  assign N3 = N13;
  assign branch_pc_high_out = (N4)? pc_r_o[21:11] : 
                              (N48)? { N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19 } : 
                              (N17)? { N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33 } : 1'b0;
  assign N4 = sel_pc;
  assign jal_pc_high_out = (N4)? pc_r_o[21:19] : 
                           (N48)? { N32, N31, N30 } : 
                           (N17)? { N46, N45, N44 } : 1'b0;
  assign pred_or_jump_addr_o = (N5)? { jal_pc_high_out, instr_o[31:31], instr_o[19:12], instr_o[20:20], instr_o[30:22] } : 
                               (N51)? jalr_prediction_i : 
                               (N50)? { branch_pc_high_out, instr_o[31:31], instr_o[7:7], instr_o[30:25], instr_o[11:9] } : 1'b0;
  assign N5 = N72;
  assign N6 = v_i & w_i;
  assign N7 = ~N6;
  assign write_branch_instr = ~N80;
  assign N80 = N78 | N79;
  assign N78 = N77 | w_instr_i[2];
  assign N77 = N76 | w_instr_i[3];
  assign N76 = N75 | w_instr_i[4];
  assign N75 = N73 | N74;
  assign N73 = ~w_instr_i[6];
  assign N74 = ~w_instr_i[5];
  assign N79 = ~w_instr_i[1];
  assign write_jal_instr = ~N92;
  assign N92 = N90 | N91;
  assign N90 = N88 | N89;
  assign N88 = N86 | N87;
  assign N86 = N84 | N85;
  assign N84 = N83 | w_instr_i[4];
  assign N83 = N81 | N82;
  assign N81 = ~w_instr_i[6];
  assign N82 = ~w_instr_i[5];
  assign N85 = ~w_instr_i[3];
  assign N87 = ~w_instr_i[2];
  assign N89 = ~w_instr_i[1];
  assign N91 = ~w_instr_i[0];
  assign N8 = write_jal_instr | write_branch_instr;
  assign N9 = ~N8;
  assign N10 = ~write_branch_instr;
  assign N11 = write_jal_instr & N10;
  assign N12 = ~write_branch_instr;
  assign N13 = v_i & N93;
  assign N93 = ~w_i;
  assign N14 = ~N13;
  assign sel_pc = ~N94;
  assign N94 = icache_data_lo_lower_sign_ ^ icache_data_lo_lower_cout_;
  assign sel_pc_p1 = N95 & icache_data_lo_lower_cout_;
  assign N95 = ~icache_data_lo_lower_sign_;
  assign N16 = sel_pc_p1 | sel_pc;
  assign N17 = ~N16;
  assign N18 = N48;
  assign N47 = ~sel_pc;
  assign N48 = sel_pc_p1 & N47;
  assign N49 = N64 | N72;
  assign N50 = ~N49;
  assign N51 = N64 & N71;

  always @(posedge clk_i) begin
    if(N52) begin
      icache_flush_r_o_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      icache_flush_r_o_sv2v_reg <= flush_i;
    end 
    if(reset_i) begin
      pc_r_o_21_sv2v_reg <= 1'b0;
      pc_r_o_20_sv2v_reg <= 1'b0;
      pc_r_o_19_sv2v_reg <= 1'b0;
      pc_r_o_18_sv2v_reg <= 1'b0;
      pc_r_o_17_sv2v_reg <= 1'b0;
      pc_r_o_16_sv2v_reg <= 1'b0;
      pc_r_o_15_sv2v_reg <= 1'b0;
      pc_r_o_14_sv2v_reg <= 1'b0;
      pc_r_o_13_sv2v_reg <= 1'b0;
      pc_r_o_12_sv2v_reg <= 1'b0;
      pc_r_o_11_sv2v_reg <= 1'b0;
      pc_r_o_10_sv2v_reg <= 1'b0;
      pc_r_o_9_sv2v_reg <= 1'b0;
      pc_r_o_8_sv2v_reg <= 1'b0;
      pc_r_o_7_sv2v_reg <= 1'b0;
      pc_r_o_6_sv2v_reg <= 1'b0;
      pc_r_o_5_sv2v_reg <= 1'b0;
      pc_r_o_4_sv2v_reg <= 1'b0;
      pc_r_o_3_sv2v_reg <= 1'b0;
      pc_r_o_2_sv2v_reg <= 1'b0;
      pc_r_o_1_sv2v_reg <= 1'b0;
      pc_r_o_0_sv2v_reg <= 1'b0;
    end else if(N15) begin
      pc_r_o_21_sv2v_reg <= pc_i[21];
      pc_r_o_20_sv2v_reg <= pc_i[20];
      pc_r_o_19_sv2v_reg <= pc_i[19];
      pc_r_o_18_sv2v_reg <= pc_i[18];
      pc_r_o_17_sv2v_reg <= pc_i[17];
      pc_r_o_16_sv2v_reg <= pc_i[16];
      pc_r_o_15_sv2v_reg <= pc_i[15];
      pc_r_o_14_sv2v_reg <= pc_i[14];
      pc_r_o_13_sv2v_reg <= pc_i[13];
      pc_r_o_12_sv2v_reg <= pc_i[12];
      pc_r_o_11_sv2v_reg <= pc_i[11];
      pc_r_o_10_sv2v_reg <= pc_i[10];
      pc_r_o_9_sv2v_reg <= pc_i[9];
      pc_r_o_8_sv2v_reg <= pc_i[8];
      pc_r_o_7_sv2v_reg <= pc_i[7];
      pc_r_o_6_sv2v_reg <= pc_i[6];
      pc_r_o_5_sv2v_reg <= pc_i[5];
      pc_r_o_4_sv2v_reg <= pc_i[4];
      pc_r_o_3_sv2v_reg <= pc_i[3];
      pc_r_o_2_sv2v_reg <= pc_i[2];
      pc_r_o_1_sv2v_reg <= pc_i[1];
      pc_r_o_0_sv2v_reg <= pc_i[0];
    end 
  end


endmodule



module cl_decode
(
  instruction_i,
  decode_o,
  fp_decode_o
);

  input [31:0] instruction_i;
  output [30:0] decode_o;
  output [10:0] fp_decode_o;
  wire [30:0] decode_o;
  wire [10:0] fp_decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,decode_o_is_amo_aq_,decode_o_is_amo_rl_,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,
  N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,
  N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,
  N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,
  N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,
  N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
  N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,
  N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,
  N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,
  N558,N559,N560,N561,N562,N563,N564,N566,N567,N568,N569,N571,N572,N573,N574,N575,
  N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,
  N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883;
  assign decode_o_is_amo_aq_ = instruction_i[26];
  assign decode_o[11] = decode_o_is_amo_aq_;
  assign decode_o_is_amo_rl_ = instruction_i[25];
  assign decode_o[10] = decode_o_is_amo_rl_;
  assign N69 = N115 | N556;
  assign N70 = N117 | N556;
  assign N71 = N100 | N461;
  assign N72 = N71 | N556;
  assign N73 = N102 | N556;
  assign N74 = N553 & N554;
  assign N75 = N74 & N456;
  assign N76 = N75 & N556;
  assign N77 = N115 | instruction_i[2];
  assign N78 = N117 | instruction_i[2];
  assign N79 = N119 | N556;
  assign N81 = N123 | instruction_i[2];
  assign N83 = N129 | instruction_i[2];
  assign N85 = instruction_i[6] & instruction_i[4];
  assign N86 = N85 & instruction_i[2];
  assign N87 = N553 & N572;
  assign N88 = N555 & instruction_i[2];
  assign N89 = N87 & N88;
  assign N90 = N554 & N572;
  assign N91 = N90 & instruction_i[2];
  assign N92 = instruction_i[5] & N572;
  assign N93 = N92 & N556;
  assign N94 = instruction_i[6] & N572;
  assign N95 = N94 & N556;
  assign N100 = N553 | N554;
  assign N101 = N556 | N558;
  assign N102 = N100 | N458;
  assign N103 = N102 | N101;
  assign N104 = instruction_i[6] & instruction_i[5];
  assign N105 = N104 & N456;
  assign N106 = N105 & N556;
  assign N107 = instruction_i[6] | instruction_i[5];
  assign N108 = instruction_i[2] | N558;
  assign N109 = N107 | N458;
  assign N110 = N109 | N108;
  assign N111 = instruction_i[6] | N554;
  assign N112 = N111 | N458;
  assign N113 = N112 | N108;
  assign N114 = N572 | instruction_i[3];
  assign N115 = N111 | N114;
  assign N116 = N115 | N108;
  assign N117 = N107 | N114;
  assign N118 = N117 | N108;
  assign N119 = N111 | N461;
  assign N120 = N119 | N101;
  assign N122 = N553 | instruction_i[5];
  assign N123 = N122 | N114;
  assign N124 = N123 | N108;
  assign N126 = N109 | N101;
  assign N127 = N112 | N101;
  assign N129 = N100 | N114;
  assign N130 = N129 | N108;
  assign N132 = instruction_i[4] & instruction_i[2];
  assign N133 = instruction_i[2] & N558;
  assign N134 = instruction_i[6] & instruction_i[3];
  assign N135 = N554 & instruction_i[3];
  assign N136 = instruction_i[6] & N554;
  assign N137 = N136 & instruction_i[2];
  assign N138 = instruction_i[3] & N556;
  assign N139 = instruction_i[4] & N558;
  assign N140 = N553 & N558;
  assign N141 = N136 & N572;
  assign N142 = N554 & N558;
  assign N146 = instruction_i[13] | N630;
  assign N147 = N747 | instruction_i[12];
  assign N151 = instruction_i[5] & instruction_i[1];
  assign N153 = N94 & N399;
  assign N154 = instruction_i[3] | instruction_i[2];
  assign N155 = N161 | N154;
  assign N156 = N155 | N558;
  assign N157 = instruction_i[6] | N572;
  assign N158 = N157 | N154;
  assign N159 = N158 | N558;
  assign N161 = instruction_i[6] | instruction_i[4];
  assign N162 = N555 | N556;
  assign N163 = N161 | N162;
  assign N164 = N163 | N558;
  assign N170 = instruction_i[14] | instruction_i[13];
  assign N171 = N170 | N630;
  assign N172 = instruction_i[14] | N747;
  assign N173 = N172 | instruction_i[12];
  assign N174 = N172 | N630;
  assign N175 = N145 | instruction_i[13];
  assign N176 = N175 | N630;
  assign N177 = N145 | N747;
  assign N178 = N177 | instruction_i[12];
  assign N179 = instruction_i[14] & instruction_i[13];
  assign N180 = N179 & instruction_i[12];
  assign N183 = N734 & N182;
  assign N184 = decode_o_is_amo_rl_ & instruction_i[14];
  assign N185 = N553 & instruction_i[5];
  assign N186 = N556 & instruction_i[1];
  assign N187 = N183 & N184;
  assign N188 = N185 & N411;
  assign N189 = N186 & instruction_i[0];
  assign N190 = N400 & N187;
  assign N191 = N188 & N189;
  assign N192 = N190 & N191;
  assign N194 = N747 & N630;
  assign N195 = N747 & instruction_i[12];
  assign N196 = instruction_i[13] & N630;
  assign N197 = instruction_i[13] & instruction_i[12];
  assign N200 = N633 & N643;
  assign N201 = N635 & N145;
  assign N202 = N572 & instruction_i[3];
  assign N203 = instruction_i[2] & instruction_i[1];
  assign N204 = N200 & N201;
  assign N205 = N196 & N185;
  assign N206 = N202 & N203;
  assign N207 = N204 & N205;
  assign N208 = N206 & instruction_i[0];
  assign N209 = N207 & N208;
  assign N211 = instruction_i[30] | N734;
  assign N213 = N634 | instruction_i[27];
  assign N215 = N634 & N734;
  assign N216 = instruction_i[30] & instruction_i[27];
  assign N220 = instruction_i[1] & instruction_i[0];
  assign N222 = N734 & N182;
  assign N223 = N799 & instruction_i[6];
  assign N224 = N222 & N223;
  assign N225 = N400 & N224;
  assign N226 = N225 & N364;
  assign N227 = instruction_i[27] & N182;
  assign N228 = N799 & instruction_i[6];
  assign N229 = N227 & N228;
  assign N230 = N400 & N229;
  assign N231 = N230 & N364;
  assign N232 = N734 & N182;
  assign N233 = N799 & instruction_i[6];
  assign N234 = N232 & N233;
  assign N235 = N407 & N234;
  assign N236 = N235 & N364;
  assign N237 = N734 & N182;
  assign N238 = N799 & N145;
  assign N239 = N237 & N238;
  assign N240 = N412 & N239;
  assign N241 = N240 & N282;
  assign N242 = N734 & N182;
  assign N243 = N799 & N145;
  assign N244 = N242 & N243;
  assign N245 = N412 & N244;
  assign N246 = N245 & N275;
  assign N247 = N734 & N182;
  assign N248 = N799 & N145;
  assign N249 = N247 & N248;
  assign N250 = N412 & N249;
  assign N251 = N250 & N268;
  assign N252 = instruction_i[27] & N182;
  assign N253 = N799 & N145;
  assign N254 = N252 & N253;
  assign N255 = N412 & N254;
  assign N256 = N255 & N282;
  assign N257 = instruction_i[27] & N182;
  assign N258 = N799 & N145;
  assign N259 = N257 & N258;
  assign N260 = N412 & N259;
  assign N261 = N260 & N275;
  assign N263 = N734 & N182;
  assign N264 = N799 & N145;
  assign N265 = N263 & N264;
  assign N266 = N196 & N136;
  assign N267 = N472 & N265;
  assign N268 = N266 & N414;
  assign N269 = N267 & N268;
  assign N270 = N734 & N182;
  assign N271 = N799 & N145;
  assign N272 = N270 & N271;
  assign N273 = N195 & N136;
  assign N274 = N472 & N272;
  assign N275 = N273 & N414;
  assign N276 = N274 & N275;
  assign N277 = N734 & N182;
  assign N278 = N799 & N145;
  assign N279 = N277 & N278;
  assign N280 = N194 & N136;
  assign N281 = N472 & N279;
  assign N282 = N280 & N414;
  assign N283 = N281 & N282;
  assign N285 = N734 & N182;
  assign N286 = N799 & N430;
  assign N287 = instruction_i[12] & instruction_i[6];
  assign N288 = N285 & N286;
  assign N289 = N448 & N287;
  assign N290 = N483 & N288;
  assign N291 = N370 & N289;
  assign N292 = N290 & N291;
  assign N293 = N292 & N364;
  assign N294 = N734 & N182;
  assign N295 = N799 & N430;
  assign N296 = N294 & N295;
  assign N297 = N438 & N296;
  assign N298 = N297 & N373;
  assign N299 = N298 & N556;
  assign N300 = N734 & N182;
  assign N301 = N799 & N430;
  assign N302 = N300 & N301;
  assign N303 = N438 & N302;
  assign N304 = N303 & N318;
  assign N305 = N304 & N556;
  assign N307 = N734 & N182;
  assign N308 = N799 & N430;
  assign N309 = N307 & N308;
  assign N310 = N479 & N309;
  assign N311 = N310 & N373;
  assign N312 = N311 & N556;
  assign N313 = N734 & N182;
  assign N314 = N799 & N430;
  assign N315 = N313 & N314;
  assign N316 = N436 & N444;
  assign N317 = N479 & N315;
  assign N318 = N316 & N371;
  assign N319 = N317 & N318;
  assign N320 = N319 & N556;
  assign N322 = N734 & N182;
  assign N323 = N799 & N430;
  assign N324 = N322 & N323;
  assign N325 = N483 & N324;
  assign N326 = N325 & N334;
  assign N327 = N326 & N364;
  assign N328 = N734 & N182;
  assign N329 = N799 & N430;
  assign N330 = N630 & instruction_i[6];
  assign N331 = N328 & N329;
  assign N332 = N448 & N330;
  assign N333 = N450 & N331;
  assign N334 = N370 & N332;
  assign N335 = N333 & N334;
  assign N336 = N335 & N364;
  assign N337 = N90 & N88;
  assign N338 = N341 & N337;
  assign N339 = N145 & instruction_i[13];
  assign N340 = N630 & N553;
  assign N341 = N339 & N340;
  assign N342 = N92 & N88;
  assign N343 = N341 & N342;
  assign N344 = N182 & N799;
  assign N345 = N344 & N136;
  assign N346 = N345 & N457;
  assign N347 = N182 & N799;
  assign N348 = N347 & N136;
  assign N349 = N456 & instruction_i[2];
  assign N350 = N348 & N349;
  assign N351 = N182 & N799;
  assign N352 = N351 & N136;
  assign N353 = N202 & N556;
  assign N354 = N352 & N353;
  assign N355 = N182 & N799;
  assign N356 = N355 & N136;
  assign N357 = N202 & instruction_i[2];
  assign N358 = N356 & N357;
  assign N360 = instruction_i[27] & N182;
  assign N361 = N799 & instruction_i[6];
  assign N362 = N554 & instruction_i[4];
  assign N363 = N360 & N361;
  assign N364 = N362 & N399;
  assign N365 = N407 & N363;
  assign N366 = N365 & N364;
  assign N367 = instruction_i[27] & N182;
  assign N368 = N799 & N430;
  assign N369 = N367 & N368;
  assign N370 = N436 & N437;
  assign N371 = N136 & N411;
  assign N372 = N468 & N369;
  assign N373 = N370 & N371;
  assign N374 = N372 & N373;
  assign N375 = N374 & N556;
  assign N392 = N182 & N799;
  assign N393 = N392 & N136;
  assign N394 = N393 & N220;
  assign N396 = N633 & N634;
  assign N397 = N643 & N635;
  assign N398 = N734 & instruction_i[4];
  assign N399 = N555 & N556;
  assign N400 = N396 & N397;
  assign N401 = N398 & N399;
  assign N402 = N400 & N401;
  assign N403 = instruction_i[27] & instruction_i[4];
  assign N404 = N403 & N399;
  assign N405 = N400 & N404;
  assign N406 = N643 & instruction_i[28];
  assign N407 = N396 & N406;
  assign N408 = N407 & N401;
  assign N409 = instruction_i[29] & N635;
  assign N410 = N734 & N145;
  assign N411 = instruction_i[4] & N555;
  assign N412 = N396 & N409;
  assign N413 = N410 & N194;
  assign N414 = N411 & N556;
  assign N415 = N412 & N413;
  assign N416 = N415 & N414;
  assign N417 = N410 & N195;
  assign N418 = N412 & N417;
  assign N419 = N418 & N414;
  assign N420 = N410 & N196;
  assign N421 = N412 & N420;
  assign N422 = N421 & N414;
  assign N423 = instruction_i[27] & N145;
  assign N424 = N423 & N194;
  assign N425 = N412 & N424;
  assign N426 = N425 & N414;
  assign N427 = N423 & N195;
  assign N428 = N412 & N427;
  assign N429 = N428 & N414;
  assign N434 = instruction_i[31] & instruction_i[30];
  assign N435 = N734 & N430;
  assign N436 = N431 & N432;
  assign N437 = N571 & N433;
  assign N438 = N434 & N406;
  assign N439 = N435 & N436;
  assign N440 = N437 & N411;
  assign N441 = N438 & N439;
  assign N442 = N440 & N556;
  assign N443 = N441 & N442;
  assign N444 = N571 & instruction_i[20];
  assign N445 = N444 & N411;
  assign N446 = N445 & N556;
  assign N447 = N441 & N446;
  assign N448 = N145 & N747;
  assign N449 = N630 & instruction_i[4];
  assign N450 = N434 & N497;
  assign N451 = N437 & N448;
  assign N452 = N449 & N399;
  assign N453 = N450 & N439;
  assign N454 = N451 & N452;
  assign N455 = N453 & N454;
  assign N456 = N572 & N555;
  assign N457 = N456 & N556;
  assign N458 = instruction_i[4] | instruction_i[3];
  assign N459 = N458 | N556;
  assign N461 = instruction_i[4] | N555;
  assign N462 = N461 | instruction_i[2];
  assign N464 = N461 | N556;
  assign N466 = N407 & N404;
  assign N467 = instruction_i[27] & N430;
  assign N468 = N522 & N406;
  assign N469 = N467 & N436;
  assign N470 = N468 & N469;
  assign N471 = N470 & N442;
  assign N472 = N500 & N409;
  assign N473 = N472 & N420;
  assign N474 = N473 & N414;
  assign N475 = N472 & N413;
  assign N476 = N475 & N414;
  assign N477 = N472 & N417;
  assign N478 = N477 & N414;
  assign N479 = N434 & N397;
  assign N480 = N479 & N439;
  assign N481 = N480 & N442;
  assign N482 = N480 & N446;
  assign N483 = N434 & N409;
  assign N484 = N498 & N399;
  assign N485 = N483 & N439;
  assign N486 = N451 & N484;
  assign N487 = N485 & N486;
  assign N488 = N485 & N454;
  assign N489 = instruction_i[4] & instruction_i[3];
  assign N490 = instruction_i[31] & instruction_i[27];
  assign N491 = N490 & instruction_i[4];
  assign N492 = instruction_i[30] & instruction_i[29];
  assign N493 = instruction_i[20] & instruction_i[4];
  assign N494 = N492 & N493;
  assign N495 = N434 & N534;
  assign N496 = N495 & instruction_i[4];
  assign N497 = instruction_i[29] & instruction_i[28];
  assign N498 = instruction_i[12] & instruction_i[4];
  assign N499 = N497 & N498;
  assign N500 = instruction_i[31] & N634;
  assign N501 = instruction_i[28] & instruction_i[4];
  assign N502 = N500 & N501;
  assign N503 = N643 & instruction_i[4];
  assign N504 = N500 & N503;
  assign N505 = instruction_i[31] & N643;
  assign N506 = instruction_i[24] & instruction_i[4];
  assign N507 = N505 & N506;
  assign N508 = instruction_i[23] & instruction_i[4];
  assign N509 = N505 & N508;
  assign N510 = instruction_i[22] & instruction_i[4];
  assign N511 = N505 & N510;
  assign N512 = instruction_i[21] & instruction_i[4];
  assign N513 = N505 & N512;
  assign N514 = instruction_i[30] & instruction_i[24];
  assign N515 = N514 & instruction_i[4];
  assign N516 = instruction_i[30] & instruction_i[23];
  assign N517 = N516 & instruction_i[4];
  assign N518 = instruction_i[30] & instruction_i[22];
  assign N519 = N518 & instruction_i[4];
  assign N520 = instruction_i[30] & instruction_i[21];
  assign N521 = N520 & instruction_i[4];
  assign N522 = N633 & instruction_i[30];
  assign N523 = N522 & N493;
  assign N524 = N635 & instruction_i[4];
  assign N525 = N522 & N524;
  assign N526 = instruction_i[29] & instruction_i[27];
  assign N527 = instruction_i[13] & instruction_i[4];
  assign N528 = N526 & N527;
  assign N529 = N522 & N398;
  assign N530 = N633 & instruction_i[29];
  assign N531 = N530 & N501;
  assign N532 = instruction_i[29] & instruction_i[14];
  assign N533 = N532 & instruction_i[4];
  assign N534 = instruction_i[29] & instruction_i[13];
  assign N535 = N534 & N498;
  assign N546 = N734 & N182;
  assign N547 = decode_o_is_amo_rl_ & N145;
  assign N548 = N546 & N547;
  assign N549 = N400 & N548;
  assign N550 = N549 & N191;
  assign N553 = ~instruction_i[6];
  assign N554 = ~instruction_i[5];
  assign N555 = ~instruction_i[3];
  assign N556 = ~instruction_i[2];
  assign N557 = ~instruction_i[1];
  assign N558 = ~instruction_i[0];
  assign N559 = N554 | N553;
  assign N560 = instruction_i[4] | N559;
  assign N561 = N555 | N560;
  assign N562 = N556 | N561;
  assign N563 = N557 | N562;
  assign N564 = N558 | N563;
  assign decode_o[21] = ~N564;
  assign N566 = instruction_i[3] | N560;
  assign N567 = N556 | N566;
  assign N568 = N557 | N567;
  assign N569 = N558 | N568;
  assign decode_o[20] = ~N569;
  assign N571 = ~instruction_i[21];
  assign N572 = ~instruction_i[4];
  assign N573 = instruction_i[30] | instruction_i[31];
  assign N574 = N643 | N573;
  assign N575 = N635 | N574;
  assign N576 = instruction_i[27] | N575;
  assign N577 = decode_o_is_amo_aq_ | N576;
  assign N578 = decode_o_is_amo_rl_ | N577;
  assign N579 = instruction_i[24] | N578;
  assign N580 = instruction_i[23] | N579;
  assign N581 = instruction_i[22] | N580;
  assign N582 = N571 | N581;
  assign N583 = instruction_i[20] | N582;
  assign N584 = instruction_i[19] | N583;
  assign N585 = instruction_i[18] | N584;
  assign N586 = instruction_i[17] | N585;
  assign N587 = instruction_i[16] | N586;
  assign N588 = instruction_i[15] | N587;
  assign N589 = instruction_i[14] | N588;
  assign N590 = instruction_i[13] | N589;
  assign N591 = instruction_i[12] | N590;
  assign N592 = instruction_i[11] | N591;
  assign N593 = instruction_i[10] | N592;
  assign N594 = instruction_i[9] | N593;
  assign N595 = instruction_i[8] | N594;
  assign N596 = instruction_i[7] | N595;
  assign N597 = N553 | N596;
  assign N598 = N554 | N597;
  assign N599 = N572 | N598;
  assign N600 = instruction_i[3] | N599;
  assign N601 = instruction_i[2] | N600;
  assign N602 = N557 | N601;
  assign N603 = N558 | N602;
  assign decode_o[1] = ~N603;
  assign N605 = instruction_i[5] | instruction_i[6];
  assign N606 = instruction_i[4] | N605;
  assign N607 = instruction_i[3] | N606;
  assign N608 = instruction_i[2] | N607;
  assign N609 = N557 | N608;
  assign N610 = N558 | N609;
  assign N611 = ~N610;
  assign N612 = N556 | N607;
  assign N613 = N557 | N612;
  assign N614 = N558 | N613;
  assign N615 = ~N614;
  assign N616 = N554 | instruction_i[6];
  assign N617 = instruction_i[4] | N616;
  assign N618 = instruction_i[3] | N617;
  assign N619 = instruction_i[2] | N618;
  assign N620 = N557 | N619;
  assign N621 = N558 | N620;
  assign N622 = ~N621;
  assign N623 = N556 | N618;
  assign N624 = N557 | N623;
  assign N625 = N558 | N624;
  assign N626 = ~N625;
  assign N627 = instruction_i[13] | instruction_i[14];
  assign N628 = instruction_i[12] | N627;
  assign N629 = ~N628;
  assign N630 = ~instruction_i[12];
  assign N631 = N630 | N627;
  assign N632 = ~N631;
  assign N633 = ~instruction_i[31];
  assign N634 = ~instruction_i[30];
  assign N635 = ~instruction_i[28];
  assign N636 = N634 | N633;
  assign N637 = instruction_i[29] | N636;
  assign N638 = N635 | N637;
  assign N639 = instruction_i[27] | N638;
  assign N640 = decode_o_is_amo_aq_ | N639;
  assign N641 = decode_o_is_amo_rl_ | N640;
  assign N642 = ~N641;
  assign N643 = ~instruction_i[29];
  assign N644 = N643 | N636;
  assign N645 = N635 | N644;
  assign N646 = instruction_i[27] | N645;
  assign N647 = decode_o_is_amo_aq_ | N646;
  assign N648 = decode_o_is_amo_rl_ | N647;
  assign N649 = ~N648;
  assign N650 = N572 | N559;
  assign N651 = instruction_i[3] | N650;
  assign N652 = instruction_i[2] | N651;
  assign N653 = N557 | N652;
  assign N654 = N558 | N653;
  assign N655 = ~N654;
  assign N656 = instruction_i[30] | N633;
  assign N657 = N643 | N656;
  assign N658 = instruction_i[28] | N657;
  assign N659 = instruction_i[27] | N658;
  assign N660 = decode_o_is_amo_aq_ | N659;
  assign N661 = decode_o_is_amo_rl_ | N660;
  assign N662 = ~N661;
  assign N663 = instruction_i[28] | N644;
  assign N664 = instruction_i[27] | N663;
  assign N665 = decode_o_is_amo_aq_ | N664;
  assign N666 = decode_o_is_amo_rl_ | N665;
  assign N667 = ~N666;
  assign N668 = instruction_i[23] | instruction_i[24];
  assign N669 = instruction_i[22] | N668;
  assign N670 = instruction_i[21] | N669;
  assign N671 = instruction_i[20] | N670;
  assign N672 = ~N671;
  assign N673 = instruction_i[28] | N637;
  assign N674 = instruction_i[27] | N673;
  assign N675 = decode_o_is_amo_aq_ | N674;
  assign N676 = decode_o_is_amo_rl_ | N675;
  assign N677 = ~N676;
  assign N678 = instruction_i[10] | instruction_i[11];
  assign N679 = instruction_i[9] | N678;
  assign N680 = instruction_i[8] | N679;
  assign N681 = instruction_i[7] | N680;
  assign N682 = ~N681;
  assign N98 = (N0)? 1'b1 : 
               (N1)? N97 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N80;
  assign N1 = N82;
  assign N2 = N84;
  assign N3 = N96;
  assign N99 = (N4)? N98 : 
               (N221)? 1'b0 : 1'b0;
  assign N4 = N220;
  assign decode_o[28] = (N5)? 1'b0 : 
                        (N6)? N99 : 1'b0;
  assign N5 = N682;
  assign N6 = N681;
  assign N149 = (N7)? N148 : 
                (N8)? 1'b0 : 1'b0;
  assign N7 = N145;
  assign N8 = instruction_i[14];
  assign N150 = (N9)? 1'b1 : 
                (N10)? N144 : 
                (N11)? 1'b1 : 
                (N12)? N149 : 
                (N13)? 1'b0 : 1'b0;
  assign N9 = N121;
  assign N10 = N125;
  assign N11 = N128;
  assign N12 = N131;
  assign N13 = N143;
  assign decode_o[30] = (N14)? N150 : 
                        (N15)? 1'b0 : 1'b0;
  assign N14 = instruction_i[1];
  assign N15 = N557;
  assign N169 = (N16)? 1'b1 : 
                (N17)? N168 : 
                (N167)? 1'b0 : 1'b0;
  assign N16 = N160;
  assign N17 = N165;
  assign decode_o[29] = (N18)? N169 : 
                        (N152)? 1'b0 : 1'b0;
  assign N18 = N151;
  assign decode_o[2] = (N19)? N181 : 
                       (N20)? 1'b0 : 1'b0;
  assign N19 = N655;
  assign N20 = N654;
  assign { N199, N198 } = (N21)? { 1'b0, 1'b0 } : 
                          (N22)? { 1'b0, 1'b1 } : 
                          (N23)? { 1'b1, 1'b0 } : 
                          (N24)? { 1'b1, 1'b1 } : 1'b0;
  assign N21 = N194;
  assign N22 = N195;
  assign N23 = N196;
  assign N24 = N197;
  assign decode_o[17:16] = (N25)? { N199, N198 } : 
                           (N193)? { 1'b0, 1'b0 } : 1'b0;
  assign N25 = decode_o[18];
  assign { N219, N218, N217 } = (N26)? { 1'b1, 1'b0, 1'b0 } : 
                                (N27)? { 1'b1, 1'b0, 1'b1 } : 
                                (N28)? { 1'b1, 1'b1, 1'b0 } : 
                                (N29)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = N212;
  assign N27 = N214;
  assign N28 = N215;
  assign N29 = N216;
  assign { decode_o[12:12], decode_o[9:8] } = (N30)? { N219, N218, N217 } : 
                                              (N210)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = N209;
  assign { N391, N390, N389, N388 } = (N31)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                      (N32)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                      (N33)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                      (N34)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                      (N35)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                      (N36)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                      (N37)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                      (N38)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N39)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N40)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                      (N41)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                      (N387)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N31 = N262;
  assign N32 = N284;
  assign N33 = N293;
  assign N34 = N306;
  assign N35 = N321;
  assign N36 = N327;
  assign N37 = N336;
  assign N38 = N338;
  assign N39 = N343;
  assign N40 = N359;
  assign N41 = N376;
  assign decode_o[7:3] = (N4)? { N391, N390, N389, N359, N388 } : 
                         (N221)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N545, N544, N543, N542, N541, N540, N539, N538, N537 } = (N42)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N43)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N44)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N45)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N46)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N47)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N48)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N49)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N50)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N51)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N52)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N53)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N54)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N55)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N56)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N59)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N60)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                                    (N61)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                                    (N62)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                    (N63)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                                    (N64)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                                    (N65)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                                    (N66)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = N402;
  assign N43 = N405;
  assign N44 = N408;
  assign N45 = N416;
  assign N46 = N419;
  assign N47 = N422;
  assign N48 = N426;
  assign N49 = N429;
  assign N50 = N443;
  assign N51 = N447;
  assign N52 = N455;
  assign N53 = N457;
  assign N54 = N460;
  assign N55 = N463;
  assign N56 = N465;
  assign N57 = N466;
  assign N58 = N471;
  assign N59 = N474;
  assign N60 = N476;
  assign N61 = N478;
  assign N62 = N481;
  assign N63 = N482;
  assign N64 = N487;
  assign N65 = N488;
  assign N66 = N536;
  assign fp_decode_o = (N67)? { N545, N544, N466, N471, N543, N542, N541, N540, N539, N538, N537 } : 
                       (N395)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = N394;
  assign decode_o[0] = (N68)? N552 : 
                       (N551)? 1'b0 : 1'b0;
  assign N68 = N550;
  assign N80 = N694 | N695;
  assign N694 = N692 | N693;
  assign N692 = N690 | N691;
  assign N690 = N689 | N76;
  assign N689 = N687 | N688;
  assign N687 = N685 | N686;
  assign N685 = N683 | N684;
  assign N683 = ~N69;
  assign N684 = ~N70;
  assign N686 = ~N72;
  assign N688 = ~N73;
  assign N691 = ~N77;
  assign N693 = ~N78;
  assign N695 = ~N79;
  assign N82 = ~N81;
  assign N84 = ~N83;
  assign N96 = N135 | N701;
  assign N701 = N489 | N700;
  assign N700 = N86 | N699;
  assign N699 = N89 | N698;
  assign N698 = N91 | N697;
  assign N697 = N138 | N696;
  assign N696 = N93 | N95;
  assign N97 = N703 | N677;
  assign N703 = N662 | N702;
  assign N702 = N667 & N672;
  assign N121 = N713 | N714;
  assign N713 = N711 | N712;
  assign N711 = N709 | N710;
  assign N709 = N707 | N708;
  assign N707 = N705 | N706;
  assign N705 = N704 | N106;
  assign N704 = ~N103;
  assign N706 = ~N110;
  assign N708 = ~N113;
  assign N710 = ~N116;
  assign N712 = ~N118;
  assign N714 = ~N120;
  assign N125 = ~N124;
  assign N128 = N715 | N716;
  assign N715 = ~N126;
  assign N716 = ~N127;
  assign N131 = ~N130;
  assign N143 = N132 | N724;
  assign N724 = N133 | N723;
  assign N723 = N134 | N722;
  assign N722 = N135 | N721;
  assign N721 = N137 | N720;
  assign N720 = N138 | N719;
  assign N719 = N139 | N718;
  assign N718 = N140 | N717;
  assign N717 = N141 | N142;
  assign N144 = N642 | N649;
  assign N145 = ~instruction_i[14];
  assign N148 = N727 | N197;
  assign N727 = N725 | N726;
  assign N725 = ~N146;
  assign N726 = ~N147;
  assign N152 = ~N151;
  assign N160 = N729 | N730;
  assign N729 = N153 | N728;
  assign N728 = ~N156;
  assign N730 = ~N159;
  assign N165 = ~N164;
  assign N166 = N165 | N160;
  assign N167 = ~N166;
  assign N168 = N742 | N746;
  assign N742 = N736 | N741;
  assign N736 = ~N735;
  assign N735 = N733 | N734;
  assign N733 = N732 | instruction_i[28];
  assign N732 = N731 | instruction_i[29];
  assign N731 = instruction_i[31] | instruction_i[30];
  assign N734 = ~instruction_i[27];
  assign N741 = ~N740;
  assign N740 = N739 | instruction_i[27];
  assign N739 = N738 | instruction_i[28];
  assign N738 = N737 | instruction_i[29];
  assign N737 = instruction_i[31] | N634;
  assign N746 = N745 & N734;
  assign N745 = N744 & N635;
  assign N744 = N743 & N643;
  assign N743 = N633 & N634;
  assign decode_o[27] = N611 | N615;
  assign decode_o[26] = N622 | N626;
  assign decode_o[25] = N749 | N750;
  assign N749 = N611 & N748;
  assign N748 = N747 & N630;
  assign N747 = ~instruction_i[13];
  assign N750 = N622 & N629;
  assign decode_o[24] = N753 | N754;
  assign N753 = N611 & N752;
  assign N752 = ~N751;
  assign N751 = instruction_i[13] | N630;
  assign N754 = N622 & N632;
  assign decode_o[23] = N611 & N756;
  assign N756 = ~N755;
  assign N755 = N145 | instruction_i[13];
  assign decode_o[22] = ~N761;
  assign N761 = N760 | N557;
  assign N760 = N759 | instruction_i[2];
  assign N759 = N758 | instruction_i[3];
  assign N758 = N757 | instruction_i[4];
  assign N757 = N553 | N554;
  assign decode_o[15] = ~N784;
  assign N784 = N783 | N558;
  assign N783 = N782 | N557;
  assign N782 = N781 | N556;
  assign N781 = N780 | N555;
  assign N780 = N779 | instruction_i[4];
  assign N779 = N778 | instruction_i[5];
  assign N778 = N777 | instruction_i[6];
  assign N777 = N776 | instruction_i[7];
  assign N776 = N775 | instruction_i[8];
  assign N775 = N774 | instruction_i[9];
  assign N774 = N773 | instruction_i[10];
  assign N773 = N772 | instruction_i[11];
  assign N772 = N771 | instruction_i[12];
  assign N771 = N770 | instruction_i[13];
  assign N770 = N769 | instruction_i[14];
  assign N769 = N768 | instruction_i[15];
  assign N768 = N767 | instruction_i[16];
  assign N767 = N766 | instruction_i[17];
  assign N766 = N765 | instruction_i[18];
  assign N765 = N764 | instruction_i[19];
  assign N764 = N763 | instruction_i[28];
  assign N763 = N762 | instruction_i[29];
  assign N762 = instruction_i[31] | instruction_i[30];
  assign N181 = N793 | N180;
  assign N793 = N791 | N792;
  assign N791 = N789 | N790;
  assign N789 = N787 | N788;
  assign N787 = N785 | N786;
  assign N785 = ~N171;
  assign N786 = ~N173;
  assign N788 = ~N174;
  assign N790 = ~N176;
  assign N792 = ~N178;
  assign decode_o[19] = ~N810;
  assign N810 = N809 | N558;
  assign N809 = N808 | N557;
  assign N808 = N807 | instruction_i[2];
  assign N807 = N806 | instruction_i[3];
  assign N806 = N805 | N572;
  assign N805 = N804 | N554;
  assign N804 = N803 | instruction_i[6];
  assign N803 = N802 | instruction_i[12];
  assign N802 = N801 | instruction_i[13];
  assign N801 = N800 | instruction_i[14];
  assign N800 = N798 | N799;
  assign N798 = N797 | decode_o_is_amo_aq_;
  assign N797 = N796 | instruction_i[27];
  assign N796 = N795 | instruction_i[28];
  assign N795 = N794 | instruction_i[29];
  assign N794 = instruction_i[31] | instruction_i[30];
  assign N799 = ~decode_o_is_amo_rl_;
  assign N182 = ~decode_o_is_amo_aq_;
  assign decode_o[18] = N192;
  assign N193 = ~decode_o[18];
  assign decode_o[13] = ~N831;
  assign N831 = N830 | N558;
  assign N830 = N829 | N557;
  assign N829 = N828 | N556;
  assign N828 = N827 | N555;
  assign N827 = N826 | instruction_i[4];
  assign N826 = N825 | N554;
  assign N825 = N824 | instruction_i[6];
  assign N824 = N823 | instruction_i[12];
  assign N823 = N822 | N747;
  assign N822 = N821 | instruction_i[14];
  assign N821 = N820 | instruction_i[20];
  assign N820 = N819 | instruction_i[21];
  assign N819 = N818 | instruction_i[22];
  assign N818 = N817 | instruction_i[23];
  assign N817 = N816 | instruction_i[24];
  assign N816 = N815 | decode_o_is_amo_rl_;
  assign N815 = N814 | decode_o_is_amo_aq_;
  assign N814 = N813 | instruction_i[27];
  assign N813 = N812 | N635;
  assign N812 = N811 | instruction_i[29];
  assign N811 = instruction_i[31] | instruction_i[30];
  assign decode_o[14] = ~N852;
  assign N852 = N851 | N558;
  assign N851 = N850 | N557;
  assign N850 = N849 | N556;
  assign N849 = N848 | N555;
  assign N848 = N847 | instruction_i[4];
  assign N847 = N846 | N554;
  assign N846 = N845 | instruction_i[6];
  assign N845 = N844 | instruction_i[12];
  assign N844 = N843 | N747;
  assign N843 = N842 | instruction_i[14];
  assign N842 = N841 | instruction_i[20];
  assign N841 = N840 | instruction_i[21];
  assign N840 = N839 | instruction_i[22];
  assign N839 = N838 | instruction_i[23];
  assign N838 = N837 | instruction_i[24];
  assign N837 = N836 | decode_o_is_amo_rl_;
  assign N836 = N835 | N182;
  assign N835 = N834 | instruction_i[27];
  assign N834 = N833 | N635;
  assign N833 = N832 | instruction_i[29];
  assign N832 = instruction_i[31] | instruction_i[30];
  assign N210 = ~N209;
  assign N212 = ~N211;
  assign N214 = ~N213;
  assign N221 = ~N220;
  assign N262 = N858 | N261;
  assign N858 = N857 | N256;
  assign N857 = N856 | N251;
  assign N856 = N855 | N246;
  assign N855 = N854 | N241;
  assign N854 = N853 | N236;
  assign N853 = N226 | N231;
  assign N284 = N859 | N283;
  assign N859 = N269 | N276;
  assign N306 = N299 | N305;
  assign N321 = N312 | N320;
  assign N359 = N861 | N358;
  assign N861 = N860 | N354;
  assign N860 = N346 | N350;
  assign N376 = N366 | N375;
  assign N377 = N284 | N262;
  assign N378 = N293 | N377;
  assign N379 = N306 | N378;
  assign N380 = N321 | N379;
  assign N381 = N327 | N380;
  assign N382 = N336 | N381;
  assign N383 = N338 | N382;
  assign N384 = N343 | N383;
  assign N385 = N359 | N384;
  assign N386 = N376 | N385;
  assign N387 = ~N386;
  assign N395 = ~N394;
  assign N430 = ~instruction_i[24];
  assign N431 = ~instruction_i[23];
  assign N432 = ~instruction_i[22];
  assign N433 = ~instruction_i[20];
  assign N460 = ~N459;
  assign N463 = ~N462;
  assign N465 = ~N464;
  assign N536 = N489 | N882;
  assign N882 = N132 | N881;
  assign N881 = N491 | N880;
  assign N880 = N494 | N879;
  assign N879 = N496 | N878;
  assign N878 = N499 | N877;
  assign N877 = N502 | N876;
  assign N876 = N504 | N875;
  assign N875 = N507 | N874;
  assign N874 = N509 | N873;
  assign N873 = N511 | N872;
  assign N872 = N513 | N871;
  assign N871 = N515 | N870;
  assign N870 = N517 | N869;
  assign N869 = N519 | N868;
  assign N868 = N521 | N867;
  assign N867 = N523 | N866;
  assign N866 = N525 | N865;
  assign N865 = N528 | N864;
  assign N864 = N529 | N863;
  assign N863 = N531 | N862;
  assign N862 = N533 | N535;
  assign N551 = ~N550;
  assign N552 = N883 | N197;
  assign N883 = N195 | N196;

endmodule



module bsg_dff_reset_width_p140
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [139:0] data_i;
  output [139:0] data_o;
  input clk_i;
  input reset_i;
  wire [139:0] data_o;
  reg data_o_139_sv2v_reg,data_o_138_sv2v_reg,data_o_137_sv2v_reg,data_o_136_sv2v_reg,
  data_o_135_sv2v_reg,data_o_134_sv2v_reg,data_o_133_sv2v_reg,data_o_132_sv2v_reg,
  data_o_131_sv2v_reg,data_o_130_sv2v_reg,data_o_129_sv2v_reg,data_o_128_sv2v_reg,
  data_o_127_sv2v_reg,data_o_126_sv2v_reg,data_o_125_sv2v_reg,data_o_124_sv2v_reg,
  data_o_123_sv2v_reg,data_o_122_sv2v_reg,data_o_121_sv2v_reg,data_o_120_sv2v_reg,
  data_o_119_sv2v_reg,data_o_118_sv2v_reg,data_o_117_sv2v_reg,data_o_116_sv2v_reg,
  data_o_115_sv2v_reg,data_o_114_sv2v_reg,data_o_113_sv2v_reg,data_o_112_sv2v_reg,
  data_o_111_sv2v_reg,data_o_110_sv2v_reg,data_o_109_sv2v_reg,data_o_108_sv2v_reg,
  data_o_107_sv2v_reg,data_o_106_sv2v_reg,data_o_105_sv2v_reg,data_o_104_sv2v_reg,
  data_o_103_sv2v_reg,data_o_102_sv2v_reg,data_o_101_sv2v_reg,data_o_100_sv2v_reg,
  data_o_99_sv2v_reg,data_o_98_sv2v_reg,data_o_97_sv2v_reg,data_o_96_sv2v_reg,
  data_o_95_sv2v_reg,data_o_94_sv2v_reg,data_o_93_sv2v_reg,data_o_92_sv2v_reg,
  data_o_91_sv2v_reg,data_o_90_sv2v_reg,data_o_89_sv2v_reg,data_o_88_sv2v_reg,
  data_o_87_sv2v_reg,data_o_86_sv2v_reg,data_o_85_sv2v_reg,data_o_84_sv2v_reg,
  data_o_83_sv2v_reg,data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,
  data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,data_o_75_sv2v_reg,
  data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,data_o_71_sv2v_reg,
  data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,data_o_67_sv2v_reg,
  data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,
  data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,
  data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,
  data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,
  data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,
  data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,
  data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,
  data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,
  data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,
  data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_139_sv2v_reg <= 1'b0;
      data_o_138_sv2v_reg <= 1'b0;
      data_o_137_sv2v_reg <= 1'b0;
      data_o_136_sv2v_reg <= 1'b0;
      data_o_135_sv2v_reg <= 1'b0;
      data_o_134_sv2v_reg <= 1'b0;
      data_o_133_sv2v_reg <= 1'b0;
      data_o_132_sv2v_reg <= 1'b0;
      data_o_131_sv2v_reg <= 1'b0;
      data_o_130_sv2v_reg <= 1'b0;
      data_o_129_sv2v_reg <= 1'b0;
      data_o_128_sv2v_reg <= 1'b0;
      data_o_127_sv2v_reg <= 1'b0;
      data_o_126_sv2v_reg <= 1'b0;
      data_o_125_sv2v_reg <= 1'b0;
      data_o_124_sv2v_reg <= 1'b0;
      data_o_123_sv2v_reg <= 1'b0;
      data_o_122_sv2v_reg <= 1'b0;
      data_o_121_sv2v_reg <= 1'b0;
      data_o_120_sv2v_reg <= 1'b0;
      data_o_119_sv2v_reg <= 1'b0;
      data_o_118_sv2v_reg <= 1'b0;
      data_o_117_sv2v_reg <= 1'b0;
      data_o_116_sv2v_reg <= 1'b0;
      data_o_115_sv2v_reg <= 1'b0;
      data_o_114_sv2v_reg <= 1'b0;
      data_o_113_sv2v_reg <= 1'b0;
      data_o_112_sv2v_reg <= 1'b0;
      data_o_111_sv2v_reg <= 1'b0;
      data_o_110_sv2v_reg <= 1'b0;
      data_o_109_sv2v_reg <= 1'b0;
      data_o_108_sv2v_reg <= 1'b0;
      data_o_107_sv2v_reg <= 1'b0;
      data_o_106_sv2v_reg <= 1'b0;
      data_o_105_sv2v_reg <= 1'b0;
      data_o_104_sv2v_reg <= 1'b0;
      data_o_103_sv2v_reg <= 1'b0;
      data_o_102_sv2v_reg <= 1'b0;
      data_o_101_sv2v_reg <= 1'b0;
      data_o_100_sv2v_reg <= 1'b0;
      data_o_99_sv2v_reg <= 1'b0;
      data_o_98_sv2v_reg <= 1'b0;
      data_o_97_sv2v_reg <= 1'b0;
      data_o_96_sv2v_reg <= 1'b0;
      data_o_95_sv2v_reg <= 1'b0;
      data_o_94_sv2v_reg <= 1'b0;
      data_o_93_sv2v_reg <= 1'b0;
      data_o_92_sv2v_reg <= 1'b0;
      data_o_91_sv2v_reg <= 1'b0;
      data_o_90_sv2v_reg <= 1'b0;
      data_o_89_sv2v_reg <= 1'b0;
      data_o_88_sv2v_reg <= 1'b0;
      data_o_87_sv2v_reg <= 1'b0;
      data_o_86_sv2v_reg <= 1'b0;
      data_o_85_sv2v_reg <= 1'b0;
      data_o_84_sv2v_reg <= 1'b0;
      data_o_83_sv2v_reg <= 1'b0;
      data_o_82_sv2v_reg <= 1'b0;
      data_o_81_sv2v_reg <= 1'b0;
      data_o_80_sv2v_reg <= 1'b0;
      data_o_79_sv2v_reg <= 1'b0;
      data_o_78_sv2v_reg <= 1'b0;
      data_o_77_sv2v_reg <= 1'b0;
      data_o_76_sv2v_reg <= 1'b0;
      data_o_75_sv2v_reg <= 1'b0;
      data_o_74_sv2v_reg <= 1'b0;
      data_o_73_sv2v_reg <= 1'b0;
      data_o_72_sv2v_reg <= 1'b0;
      data_o_71_sv2v_reg <= 1'b0;
      data_o_70_sv2v_reg <= 1'b0;
      data_o_69_sv2v_reg <= 1'b0;
      data_o_68_sv2v_reg <= 1'b0;
      data_o_67_sv2v_reg <= 1'b0;
      data_o_66_sv2v_reg <= 1'b0;
      data_o_65_sv2v_reg <= 1'b0;
      data_o_64_sv2v_reg <= 1'b0;
      data_o_63_sv2v_reg <= 1'b0;
      data_o_62_sv2v_reg <= 1'b0;
      data_o_61_sv2v_reg <= 1'b0;
      data_o_60_sv2v_reg <= 1'b0;
      data_o_59_sv2v_reg <= 1'b0;
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module regfile_synth_width_p32_els_p32_num_rs_p2_x0_tied_to_zero_p1
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [4:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_v_i;
  input [9:0] r_addr_i;
  output [63:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  wire [63:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,\xz.mem_with_zero_31__31_ ,
  \xz.mem_with_zero_31__30_ ,\xz.mem_with_zero_31__29_ ,\xz.mem_with_zero_31__28_ ,
  \xz.mem_with_zero_31__27_ ,\xz.mem_with_zero_31__26_ ,\xz.mem_with_zero_31__25_ ,
  \xz.mem_with_zero_31__24_ ,\xz.mem_with_zero_31__23_ ,\xz.mem_with_zero_31__22_ ,
  \xz.mem_with_zero_31__21_ ,\xz.mem_with_zero_31__20_ ,\xz.mem_with_zero_31__19_ ,
  \xz.mem_with_zero_31__18_ ,\xz.mem_with_zero_31__17_ ,\xz.mem_with_zero_31__16_ ,
  \xz.mem_with_zero_31__15_ ,\xz.mem_with_zero_31__14_ ,\xz.mem_with_zero_31__13_ ,
  \xz.mem_with_zero_31__12_ ,\xz.mem_with_zero_31__11_ ,\xz.mem_with_zero_31__10_ ,
  \xz.mem_with_zero_31__9_ ,\xz.mem_with_zero_31__8_ ,\xz.mem_with_zero_31__7_ ,
  \xz.mem_with_zero_31__6_ ,\xz.mem_with_zero_31__5_ ,\xz.mem_with_zero_31__4_ ,
  \xz.mem_with_zero_31__3_ ,\xz.mem_with_zero_31__2_ ,\xz.mem_with_zero_31__1_ ,
  \xz.mem_with_zero_31__0_ ,\xz.mem_with_zero_30__31_ ,\xz.mem_with_zero_30__30_ ,
  \xz.mem_with_zero_30__29_ ,\xz.mem_with_zero_30__28_ ,\xz.mem_with_zero_30__27_ ,
  \xz.mem_with_zero_30__26_ ,\xz.mem_with_zero_30__25_ ,\xz.mem_with_zero_30__24_ ,
  \xz.mem_with_zero_30__23_ ,\xz.mem_with_zero_30__22_ ,\xz.mem_with_zero_30__21_ ,
  \xz.mem_with_zero_30__20_ ,\xz.mem_with_zero_30__19_ ,\xz.mem_with_zero_30__18_ ,
  \xz.mem_with_zero_30__17_ ,\xz.mem_with_zero_30__16_ ,\xz.mem_with_zero_30__15_ ,
  \xz.mem_with_zero_30__14_ ,\xz.mem_with_zero_30__13_ ,\xz.mem_with_zero_30__12_ ,
  \xz.mem_with_zero_30__11_ ,\xz.mem_with_zero_30__10_ ,\xz.mem_with_zero_30__9_ ,
  \xz.mem_with_zero_30__8_ ,\xz.mem_with_zero_30__7_ ,\xz.mem_with_zero_30__6_ ,
  \xz.mem_with_zero_30__5_ ,\xz.mem_with_zero_30__4_ ,\xz.mem_with_zero_30__3_ ,
  \xz.mem_with_zero_30__2_ ,\xz.mem_with_zero_30__1_ ,\xz.mem_with_zero_30__0_ ,
  \xz.mem_with_zero_29__31_ ,\xz.mem_with_zero_29__30_ ,\xz.mem_with_zero_29__29_ ,
  \xz.mem_with_zero_29__28_ ,\xz.mem_with_zero_29__27_ ,\xz.mem_with_zero_29__26_ ,
  \xz.mem_with_zero_29__25_ ,\xz.mem_with_zero_29__24_ ,\xz.mem_with_zero_29__23_ ,
  \xz.mem_with_zero_29__22_ ,\xz.mem_with_zero_29__21_ ,\xz.mem_with_zero_29__20_ ,
  \xz.mem_with_zero_29__19_ ,\xz.mem_with_zero_29__18_ ,\xz.mem_with_zero_29__17_ ,
  \xz.mem_with_zero_29__16_ ,\xz.mem_with_zero_29__15_ ,\xz.mem_with_zero_29__14_ ,
  \xz.mem_with_zero_29__13_ ,\xz.mem_with_zero_29__12_ ,\xz.mem_with_zero_29__11_ ,
  \xz.mem_with_zero_29__10_ ,\xz.mem_with_zero_29__9_ ,\xz.mem_with_zero_29__8_ ,
  \xz.mem_with_zero_29__7_ ,\xz.mem_with_zero_29__6_ ,\xz.mem_with_zero_29__5_ ,
  \xz.mem_with_zero_29__4_ ,\xz.mem_with_zero_29__3_ ,\xz.mem_with_zero_29__2_ ,
  \xz.mem_with_zero_29__1_ ,\xz.mem_with_zero_29__0_ ,\xz.mem_with_zero_28__31_ ,
  \xz.mem_with_zero_28__30_ ,\xz.mem_with_zero_28__29_ ,\xz.mem_with_zero_28__28_ ,
  \xz.mem_with_zero_28__27_ ,\xz.mem_with_zero_28__26_ ,\xz.mem_with_zero_28__25_ ,
  \xz.mem_with_zero_28__24_ ,\xz.mem_with_zero_28__23_ ,\xz.mem_with_zero_28__22_ ,
  \xz.mem_with_zero_28__21_ ,\xz.mem_with_zero_28__20_ ,\xz.mem_with_zero_28__19_ ,
  \xz.mem_with_zero_28__18_ ,\xz.mem_with_zero_28__17_ ,\xz.mem_with_zero_28__16_ ,
  \xz.mem_with_zero_28__15_ ,\xz.mem_with_zero_28__14_ ,\xz.mem_with_zero_28__13_ ,
  \xz.mem_with_zero_28__12_ ,\xz.mem_with_zero_28__11_ ,\xz.mem_with_zero_28__10_ ,
  \xz.mem_with_zero_28__9_ ,\xz.mem_with_zero_28__8_ ,\xz.mem_with_zero_28__7_ ,
  \xz.mem_with_zero_28__6_ ,\xz.mem_with_zero_28__5_ ,\xz.mem_with_zero_28__4_ ,
  \xz.mem_with_zero_28__3_ ,\xz.mem_with_zero_28__2_ ,\xz.mem_with_zero_28__1_ ,
  \xz.mem_with_zero_28__0_ ,\xz.mem_with_zero_27__31_ ,\xz.mem_with_zero_27__30_ ,
  \xz.mem_with_zero_27__29_ ,\xz.mem_with_zero_27__28_ ,\xz.mem_with_zero_27__27_ ,
  \xz.mem_with_zero_27__26_ ,\xz.mem_with_zero_27__25_ ,\xz.mem_with_zero_27__24_ ,
  \xz.mem_with_zero_27__23_ ,\xz.mem_with_zero_27__22_ ,\xz.mem_with_zero_27__21_ ,
  \xz.mem_with_zero_27__20_ ,\xz.mem_with_zero_27__19_ ,\xz.mem_with_zero_27__18_ ,
  \xz.mem_with_zero_27__17_ ,\xz.mem_with_zero_27__16_ ,\xz.mem_with_zero_27__15_ ,
  \xz.mem_with_zero_27__14_ ,\xz.mem_with_zero_27__13_ ,\xz.mem_with_zero_27__12_ ,
  \xz.mem_with_zero_27__11_ ,\xz.mem_with_zero_27__10_ ,\xz.mem_with_zero_27__9_ ,
  \xz.mem_with_zero_27__8_ ,\xz.mem_with_zero_27__7_ ,\xz.mem_with_zero_27__6_ ,
  \xz.mem_with_zero_27__5_ ,\xz.mem_with_zero_27__4_ ,\xz.mem_with_zero_27__3_ ,
  \xz.mem_with_zero_27__2_ ,\xz.mem_with_zero_27__1_ ,\xz.mem_with_zero_27__0_ ,
  \xz.mem_with_zero_26__31_ ,\xz.mem_with_zero_26__30_ ,\xz.mem_with_zero_26__29_ ,
  \xz.mem_with_zero_26__28_ ,\xz.mem_with_zero_26__27_ ,\xz.mem_with_zero_26__26_ ,
  \xz.mem_with_zero_26__25_ ,\xz.mem_with_zero_26__24_ ,\xz.mem_with_zero_26__23_ ,
  \xz.mem_with_zero_26__22_ ,\xz.mem_with_zero_26__21_ ,\xz.mem_with_zero_26__20_ ,
  \xz.mem_with_zero_26__19_ ,\xz.mem_with_zero_26__18_ ,\xz.mem_with_zero_26__17_ ,
  \xz.mem_with_zero_26__16_ ,\xz.mem_with_zero_26__15_ ,\xz.mem_with_zero_26__14_ ,
  \xz.mem_with_zero_26__13_ ,\xz.mem_with_zero_26__12_ ,\xz.mem_with_zero_26__11_ ,
  \xz.mem_with_zero_26__10_ ,\xz.mem_with_zero_26__9_ ,\xz.mem_with_zero_26__8_ ,
  \xz.mem_with_zero_26__7_ ,\xz.mem_with_zero_26__6_ ,\xz.mem_with_zero_26__5_ ,
  \xz.mem_with_zero_26__4_ ,\xz.mem_with_zero_26__3_ ,\xz.mem_with_zero_26__2_ ,
  \xz.mem_with_zero_26__1_ ,\xz.mem_with_zero_26__0_ ,\xz.mem_with_zero_25__31_ ,
  \xz.mem_with_zero_25__30_ ,\xz.mem_with_zero_25__29_ ,\xz.mem_with_zero_25__28_ ,
  \xz.mem_with_zero_25__27_ ,\xz.mem_with_zero_25__26_ ,\xz.mem_with_zero_25__25_ ,
  \xz.mem_with_zero_25__24_ ,\xz.mem_with_zero_25__23_ ,\xz.mem_with_zero_25__22_ ,
  \xz.mem_with_zero_25__21_ ,\xz.mem_with_zero_25__20_ ,\xz.mem_with_zero_25__19_ ,
  \xz.mem_with_zero_25__18_ ,\xz.mem_with_zero_25__17_ ,\xz.mem_with_zero_25__16_ ,
  \xz.mem_with_zero_25__15_ ,\xz.mem_with_zero_25__14_ ,\xz.mem_with_zero_25__13_ ,
  \xz.mem_with_zero_25__12_ ,\xz.mem_with_zero_25__11_ ,\xz.mem_with_zero_25__10_ ,
  \xz.mem_with_zero_25__9_ ,\xz.mem_with_zero_25__8_ ,\xz.mem_with_zero_25__7_ ,
  \xz.mem_with_zero_25__6_ ,\xz.mem_with_zero_25__5_ ,\xz.mem_with_zero_25__4_ ,
  \xz.mem_with_zero_25__3_ ,\xz.mem_with_zero_25__2_ ,\xz.mem_with_zero_25__1_ ,
  \xz.mem_with_zero_25__0_ ,\xz.mem_with_zero_24__31_ ,\xz.mem_with_zero_24__30_ ,
  \xz.mem_with_zero_24__29_ ,\xz.mem_with_zero_24__28_ ,\xz.mem_with_zero_24__27_ ,
  \xz.mem_with_zero_24__26_ ,\xz.mem_with_zero_24__25_ ,\xz.mem_with_zero_24__24_ ,
  \xz.mem_with_zero_24__23_ ,\xz.mem_with_zero_24__22_ ,\xz.mem_with_zero_24__21_ ,
  \xz.mem_with_zero_24__20_ ,\xz.mem_with_zero_24__19_ ,\xz.mem_with_zero_24__18_ ,
  \xz.mem_with_zero_24__17_ ,\xz.mem_with_zero_24__16_ ,\xz.mem_with_zero_24__15_ ,
  \xz.mem_with_zero_24__14_ ,\xz.mem_with_zero_24__13_ ,\xz.mem_with_zero_24__12_ ,
  \xz.mem_with_zero_24__11_ ,\xz.mem_with_zero_24__10_ ,\xz.mem_with_zero_24__9_ ,
  \xz.mem_with_zero_24__8_ ,\xz.mem_with_zero_24__7_ ,\xz.mem_with_zero_24__6_ ,
  \xz.mem_with_zero_24__5_ ,\xz.mem_with_zero_24__4_ ,\xz.mem_with_zero_24__3_ ,
  \xz.mem_with_zero_24__2_ ,\xz.mem_with_zero_24__1_ ,\xz.mem_with_zero_24__0_ ,
  \xz.mem_with_zero_23__31_ ,\xz.mem_with_zero_23__30_ ,\xz.mem_with_zero_23__29_ ,
  \xz.mem_with_zero_23__28_ ,\xz.mem_with_zero_23__27_ ,\xz.mem_with_zero_23__26_ ,
  \xz.mem_with_zero_23__25_ ,\xz.mem_with_zero_23__24_ ,\xz.mem_with_zero_23__23_ ,
  \xz.mem_with_zero_23__22_ ,\xz.mem_with_zero_23__21_ ,\xz.mem_with_zero_23__20_ ,
  \xz.mem_with_zero_23__19_ ,\xz.mem_with_zero_23__18_ ,\xz.mem_with_zero_23__17_ ,
  \xz.mem_with_zero_23__16_ ,\xz.mem_with_zero_23__15_ ,\xz.mem_with_zero_23__14_ ,
  \xz.mem_with_zero_23__13_ ,\xz.mem_with_zero_23__12_ ,\xz.mem_with_zero_23__11_ ,
  \xz.mem_with_zero_23__10_ ,\xz.mem_with_zero_23__9_ ,\xz.mem_with_zero_23__8_ ,
  \xz.mem_with_zero_23__7_ ,\xz.mem_with_zero_23__6_ ,\xz.mem_with_zero_23__5_ ,
  \xz.mem_with_zero_23__4_ ,\xz.mem_with_zero_23__3_ ,\xz.mem_with_zero_23__2_ ,
  \xz.mem_with_zero_23__1_ ,\xz.mem_with_zero_23__0_ ,\xz.mem_with_zero_22__31_ ,
  \xz.mem_with_zero_22__30_ ,\xz.mem_with_zero_22__29_ ,\xz.mem_with_zero_22__28_ ,
  \xz.mem_with_zero_22__27_ ,\xz.mem_with_zero_22__26_ ,\xz.mem_with_zero_22__25_ ,
  \xz.mem_with_zero_22__24_ ,\xz.mem_with_zero_22__23_ ,\xz.mem_with_zero_22__22_ ,
  \xz.mem_with_zero_22__21_ ,\xz.mem_with_zero_22__20_ ,\xz.mem_with_zero_22__19_ ,
  \xz.mem_with_zero_22__18_ ,\xz.mem_with_zero_22__17_ ,\xz.mem_with_zero_22__16_ ,
  \xz.mem_with_zero_22__15_ ,\xz.mem_with_zero_22__14_ ,\xz.mem_with_zero_22__13_ ,
  \xz.mem_with_zero_22__12_ ,\xz.mem_with_zero_22__11_ ,\xz.mem_with_zero_22__10_ ,
  \xz.mem_with_zero_22__9_ ,\xz.mem_with_zero_22__8_ ,\xz.mem_with_zero_22__7_ ,
  \xz.mem_with_zero_22__6_ ,\xz.mem_with_zero_22__5_ ,\xz.mem_with_zero_22__4_ ,
  \xz.mem_with_zero_22__3_ ,\xz.mem_with_zero_22__2_ ,\xz.mem_with_zero_22__1_ ,
  \xz.mem_with_zero_22__0_ ,\xz.mem_with_zero_21__31_ ,\xz.mem_with_zero_21__30_ ,
  \xz.mem_with_zero_21__29_ ,\xz.mem_with_zero_21__28_ ,\xz.mem_with_zero_21__27_ ,
  \xz.mem_with_zero_21__26_ ,\xz.mem_with_zero_21__25_ ,\xz.mem_with_zero_21__24_ ,
  \xz.mem_with_zero_21__23_ ,\xz.mem_with_zero_21__22_ ,\xz.mem_with_zero_21__21_ ,
  \xz.mem_with_zero_21__20_ ,\xz.mem_with_zero_21__19_ ,\xz.mem_with_zero_21__18_ ,
  \xz.mem_with_zero_21__17_ ,\xz.mem_with_zero_21__16_ ,\xz.mem_with_zero_21__15_ ,
  \xz.mem_with_zero_21__14_ ,\xz.mem_with_zero_21__13_ ,\xz.mem_with_zero_21__12_ ,
  \xz.mem_with_zero_21__11_ ,\xz.mem_with_zero_21__10_ ,\xz.mem_with_zero_21__9_ ,
  \xz.mem_with_zero_21__8_ ,\xz.mem_with_zero_21__7_ ,\xz.mem_with_zero_21__6_ ,
  \xz.mem_with_zero_21__5_ ,\xz.mem_with_zero_21__4_ ,\xz.mem_with_zero_21__3_ ,
  \xz.mem_with_zero_21__2_ ,\xz.mem_with_zero_21__1_ ,\xz.mem_with_zero_21__0_ ,
  \xz.mem_with_zero_20__31_ ,\xz.mem_with_zero_20__30_ ,\xz.mem_with_zero_20__29_ ,
  \xz.mem_with_zero_20__28_ ,\xz.mem_with_zero_20__27_ ,\xz.mem_with_zero_20__26_ ,
  \xz.mem_with_zero_20__25_ ,\xz.mem_with_zero_20__24_ ,\xz.mem_with_zero_20__23_ ,
  \xz.mem_with_zero_20__22_ ,\xz.mem_with_zero_20__21_ ,\xz.mem_with_zero_20__20_ ,
  \xz.mem_with_zero_20__19_ ,\xz.mem_with_zero_20__18_ ,\xz.mem_with_zero_20__17_ ,
  \xz.mem_with_zero_20__16_ ,\xz.mem_with_zero_20__15_ ,\xz.mem_with_zero_20__14_ ,
  \xz.mem_with_zero_20__13_ ,\xz.mem_with_zero_20__12_ ,\xz.mem_with_zero_20__11_ ,
  \xz.mem_with_zero_20__10_ ,\xz.mem_with_zero_20__9_ ,\xz.mem_with_zero_20__8_ ,
  \xz.mem_with_zero_20__7_ ,\xz.mem_with_zero_20__6_ ,\xz.mem_with_zero_20__5_ ,
  \xz.mem_with_zero_20__4_ ,\xz.mem_with_zero_20__3_ ,\xz.mem_with_zero_20__2_ ,
  \xz.mem_with_zero_20__1_ ,\xz.mem_with_zero_20__0_ ,\xz.mem_with_zero_19__31_ ,
  \xz.mem_with_zero_19__30_ ,\xz.mem_with_zero_19__29_ ,\xz.mem_with_zero_19__28_ ,
  \xz.mem_with_zero_19__27_ ,\xz.mem_with_zero_19__26_ ,\xz.mem_with_zero_19__25_ ,
  \xz.mem_with_zero_19__24_ ,\xz.mem_with_zero_19__23_ ,\xz.mem_with_zero_19__22_ ,
  \xz.mem_with_zero_19__21_ ,\xz.mem_with_zero_19__20_ ,\xz.mem_with_zero_19__19_ ,
  \xz.mem_with_zero_19__18_ ,\xz.mem_with_zero_19__17_ ,\xz.mem_with_zero_19__16_ ,
  \xz.mem_with_zero_19__15_ ,\xz.mem_with_zero_19__14_ ,\xz.mem_with_zero_19__13_ ,
  \xz.mem_with_zero_19__12_ ,\xz.mem_with_zero_19__11_ ,\xz.mem_with_zero_19__10_ ,
  \xz.mem_with_zero_19__9_ ,\xz.mem_with_zero_19__8_ ,\xz.mem_with_zero_19__7_ ,
  \xz.mem_with_zero_19__6_ ,\xz.mem_with_zero_19__5_ ,\xz.mem_with_zero_19__4_ ,
  \xz.mem_with_zero_19__3_ ,\xz.mem_with_zero_19__2_ ,\xz.mem_with_zero_19__1_ ,
  \xz.mem_with_zero_19__0_ ,\xz.mem_with_zero_18__31_ ,\xz.mem_with_zero_18__30_ ,
  \xz.mem_with_zero_18__29_ ,\xz.mem_with_zero_18__28_ ,\xz.mem_with_zero_18__27_ ,
  \xz.mem_with_zero_18__26_ ,\xz.mem_with_zero_18__25_ ,\xz.mem_with_zero_18__24_ ,
  \xz.mem_with_zero_18__23_ ,\xz.mem_with_zero_18__22_ ,\xz.mem_with_zero_18__21_ ,
  \xz.mem_with_zero_18__20_ ,\xz.mem_with_zero_18__19_ ,\xz.mem_with_zero_18__18_ ,
  \xz.mem_with_zero_18__17_ ,\xz.mem_with_zero_18__16_ ,\xz.mem_with_zero_18__15_ ,
  \xz.mem_with_zero_18__14_ ,\xz.mem_with_zero_18__13_ ,\xz.mem_with_zero_18__12_ ,
  \xz.mem_with_zero_18__11_ ,\xz.mem_with_zero_18__10_ ,\xz.mem_with_zero_18__9_ ,
  \xz.mem_with_zero_18__8_ ,\xz.mem_with_zero_18__7_ ,\xz.mem_with_zero_18__6_ ,
  \xz.mem_with_zero_18__5_ ,\xz.mem_with_zero_18__4_ ,\xz.mem_with_zero_18__3_ ,
  \xz.mem_with_zero_18__2_ ,\xz.mem_with_zero_18__1_ ,\xz.mem_with_zero_18__0_ ,
  \xz.mem_with_zero_17__31_ ,\xz.mem_with_zero_17__30_ ,\xz.mem_with_zero_17__29_ ,
  \xz.mem_with_zero_17__28_ ,\xz.mem_with_zero_17__27_ ,\xz.mem_with_zero_17__26_ ,
  \xz.mem_with_zero_17__25_ ,\xz.mem_with_zero_17__24_ ,\xz.mem_with_zero_17__23_ ,
  \xz.mem_with_zero_17__22_ ,\xz.mem_with_zero_17__21_ ,\xz.mem_with_zero_17__20_ ,
  \xz.mem_with_zero_17__19_ ,\xz.mem_with_zero_17__18_ ,\xz.mem_with_zero_17__17_ ,
  \xz.mem_with_zero_17__16_ ,\xz.mem_with_zero_17__15_ ,\xz.mem_with_zero_17__14_ ,
  \xz.mem_with_zero_17__13_ ,\xz.mem_with_zero_17__12_ ,\xz.mem_with_zero_17__11_ ,
  \xz.mem_with_zero_17__10_ ,\xz.mem_with_zero_17__9_ ,\xz.mem_with_zero_17__8_ ,
  \xz.mem_with_zero_17__7_ ,\xz.mem_with_zero_17__6_ ,\xz.mem_with_zero_17__5_ ,
  \xz.mem_with_zero_17__4_ ,\xz.mem_with_zero_17__3_ ,\xz.mem_with_zero_17__2_ ,
  \xz.mem_with_zero_17__1_ ,\xz.mem_with_zero_17__0_ ,\xz.mem_with_zero_16__31_ ,
  \xz.mem_with_zero_16__30_ ,\xz.mem_with_zero_16__29_ ,\xz.mem_with_zero_16__28_ ,
  \xz.mem_with_zero_16__27_ ,\xz.mem_with_zero_16__26_ ,\xz.mem_with_zero_16__25_ ,
  \xz.mem_with_zero_16__24_ ,\xz.mem_with_zero_16__23_ ,\xz.mem_with_zero_16__22_ ,
  \xz.mem_with_zero_16__21_ ,\xz.mem_with_zero_16__20_ ,\xz.mem_with_zero_16__19_ ,
  \xz.mem_with_zero_16__18_ ,\xz.mem_with_zero_16__17_ ,\xz.mem_with_zero_16__16_ ,
  \xz.mem_with_zero_16__15_ ,\xz.mem_with_zero_16__14_ ,\xz.mem_with_zero_16__13_ ,
  \xz.mem_with_zero_16__12_ ,\xz.mem_with_zero_16__11_ ,\xz.mem_with_zero_16__10_ ,
  \xz.mem_with_zero_16__9_ ,\xz.mem_with_zero_16__8_ ,\xz.mem_with_zero_16__7_ ,
  \xz.mem_with_zero_16__6_ ,\xz.mem_with_zero_16__5_ ,\xz.mem_with_zero_16__4_ ,
  \xz.mem_with_zero_16__3_ ,\xz.mem_with_zero_16__2_ ,\xz.mem_with_zero_16__1_ ,
  \xz.mem_with_zero_16__0_ ,\xz.mem_with_zero_15__31_ ,\xz.mem_with_zero_15__30_ ,
  \xz.mem_with_zero_15__29_ ,\xz.mem_with_zero_15__28_ ,\xz.mem_with_zero_15__27_ ,
  \xz.mem_with_zero_15__26_ ,\xz.mem_with_zero_15__25_ ,\xz.mem_with_zero_15__24_ ,
  \xz.mem_with_zero_15__23_ ,\xz.mem_with_zero_15__22_ ,\xz.mem_with_zero_15__21_ ,
  \xz.mem_with_zero_15__20_ ,\xz.mem_with_zero_15__19_ ,\xz.mem_with_zero_15__18_ ,
  \xz.mem_with_zero_15__17_ ,\xz.mem_with_zero_15__16_ ,\xz.mem_with_zero_15__15_ ,
  \xz.mem_with_zero_15__14_ ,\xz.mem_with_zero_15__13_ ,\xz.mem_with_zero_15__12_ ,
  \xz.mem_with_zero_15__11_ ,\xz.mem_with_zero_15__10_ ,\xz.mem_with_zero_15__9_ ,
  \xz.mem_with_zero_15__8_ ,\xz.mem_with_zero_15__7_ ,\xz.mem_with_zero_15__6_ ,
  \xz.mem_with_zero_15__5_ ,\xz.mem_with_zero_15__4_ ,\xz.mem_with_zero_15__3_ ,
  \xz.mem_with_zero_15__2_ ,\xz.mem_with_zero_15__1_ ,\xz.mem_with_zero_15__0_ ,
  \xz.mem_with_zero_14__31_ ,\xz.mem_with_zero_14__30_ ,\xz.mem_with_zero_14__29_ ,
  \xz.mem_with_zero_14__28_ ,\xz.mem_with_zero_14__27_ ,\xz.mem_with_zero_14__26_ ,
  \xz.mem_with_zero_14__25_ ,\xz.mem_with_zero_14__24_ ,\xz.mem_with_zero_14__23_ ,
  \xz.mem_with_zero_14__22_ ,\xz.mem_with_zero_14__21_ ,\xz.mem_with_zero_14__20_ ,
  \xz.mem_with_zero_14__19_ ,\xz.mem_with_zero_14__18_ ,\xz.mem_with_zero_14__17_ ,
  \xz.mem_with_zero_14__16_ ,\xz.mem_with_zero_14__15_ ,\xz.mem_with_zero_14__14_ ,
  \xz.mem_with_zero_14__13_ ,\xz.mem_with_zero_14__12_ ,\xz.mem_with_zero_14__11_ ,
  \xz.mem_with_zero_14__10_ ,\xz.mem_with_zero_14__9_ ,\xz.mem_with_zero_14__8_ ,
  \xz.mem_with_zero_14__7_ ,\xz.mem_with_zero_14__6_ ,\xz.mem_with_zero_14__5_ ,
  \xz.mem_with_zero_14__4_ ,\xz.mem_with_zero_14__3_ ,\xz.mem_with_zero_14__2_ ,
  \xz.mem_with_zero_14__1_ ,\xz.mem_with_zero_14__0_ ,\xz.mem_with_zero_13__31_ ,
  \xz.mem_with_zero_13__30_ ,\xz.mem_with_zero_13__29_ ,\xz.mem_with_zero_13__28_ ,
  \xz.mem_with_zero_13__27_ ,\xz.mem_with_zero_13__26_ ,\xz.mem_with_zero_13__25_ ,
  \xz.mem_with_zero_13__24_ ,\xz.mem_with_zero_13__23_ ,\xz.mem_with_zero_13__22_ ,
  \xz.mem_with_zero_13__21_ ,\xz.mem_with_zero_13__20_ ,\xz.mem_with_zero_13__19_ ,
  \xz.mem_with_zero_13__18_ ,\xz.mem_with_zero_13__17_ ,\xz.mem_with_zero_13__16_ ,
  \xz.mem_with_zero_13__15_ ,\xz.mem_with_zero_13__14_ ,\xz.mem_with_zero_13__13_ ,
  \xz.mem_with_zero_13__12_ ,\xz.mem_with_zero_13__11_ ,\xz.mem_with_zero_13__10_ ,
  \xz.mem_with_zero_13__9_ ,\xz.mem_with_zero_13__8_ ,\xz.mem_with_zero_13__7_ ,
  \xz.mem_with_zero_13__6_ ,\xz.mem_with_zero_13__5_ ,\xz.mem_with_zero_13__4_ ,
  \xz.mem_with_zero_13__3_ ,\xz.mem_with_zero_13__2_ ,\xz.mem_with_zero_13__1_ ,
  \xz.mem_with_zero_13__0_ ,\xz.mem_with_zero_12__31_ ,\xz.mem_with_zero_12__30_ ,
  \xz.mem_with_zero_12__29_ ,\xz.mem_with_zero_12__28_ ,\xz.mem_with_zero_12__27_ ,
  \xz.mem_with_zero_12__26_ ,\xz.mem_with_zero_12__25_ ,\xz.mem_with_zero_12__24_ ,
  \xz.mem_with_zero_12__23_ ,\xz.mem_with_zero_12__22_ ,\xz.mem_with_zero_12__21_ ,
  \xz.mem_with_zero_12__20_ ,\xz.mem_with_zero_12__19_ ,\xz.mem_with_zero_12__18_ ,
  \xz.mem_with_zero_12__17_ ,\xz.mem_with_zero_12__16_ ,\xz.mem_with_zero_12__15_ ,
  \xz.mem_with_zero_12__14_ ,\xz.mem_with_zero_12__13_ ,\xz.mem_with_zero_12__12_ ,
  \xz.mem_with_zero_12__11_ ,\xz.mem_with_zero_12__10_ ,\xz.mem_with_zero_12__9_ ,
  \xz.mem_with_zero_12__8_ ,\xz.mem_with_zero_12__7_ ,\xz.mem_with_zero_12__6_ ,
  \xz.mem_with_zero_12__5_ ,\xz.mem_with_zero_12__4_ ,\xz.mem_with_zero_12__3_ ,
  \xz.mem_with_zero_12__2_ ,\xz.mem_with_zero_12__1_ ,\xz.mem_with_zero_12__0_ ,
  \xz.mem_with_zero_11__31_ ,\xz.mem_with_zero_11__30_ ,\xz.mem_with_zero_11__29_ ,
  \xz.mem_with_zero_11__28_ ,\xz.mem_with_zero_11__27_ ,\xz.mem_with_zero_11__26_ ,
  \xz.mem_with_zero_11__25_ ,\xz.mem_with_zero_11__24_ ,\xz.mem_with_zero_11__23_ ,
  \xz.mem_with_zero_11__22_ ,\xz.mem_with_zero_11__21_ ,\xz.mem_with_zero_11__20_ ,
  \xz.mem_with_zero_11__19_ ,\xz.mem_with_zero_11__18_ ,\xz.mem_with_zero_11__17_ ,
  \xz.mem_with_zero_11__16_ ,\xz.mem_with_zero_11__15_ ,\xz.mem_with_zero_11__14_ ,
  \xz.mem_with_zero_11__13_ ,\xz.mem_with_zero_11__12_ ,\xz.mem_with_zero_11__11_ ,
  \xz.mem_with_zero_11__10_ ,\xz.mem_with_zero_11__9_ ,\xz.mem_with_zero_11__8_ ,
  \xz.mem_with_zero_11__7_ ,\xz.mem_with_zero_11__6_ ,\xz.mem_with_zero_11__5_ ,
  \xz.mem_with_zero_11__4_ ,\xz.mem_with_zero_11__3_ ,\xz.mem_with_zero_11__2_ ,
  \xz.mem_with_zero_11__1_ ,\xz.mem_with_zero_11__0_ ,\xz.mem_with_zero_10__31_ ,
  \xz.mem_with_zero_10__30_ ,\xz.mem_with_zero_10__29_ ,\xz.mem_with_zero_10__28_ ,
  \xz.mem_with_zero_10__27_ ,\xz.mem_with_zero_10__26_ ,\xz.mem_with_zero_10__25_ ,
  \xz.mem_with_zero_10__24_ ,\xz.mem_with_zero_10__23_ ,\xz.mem_with_zero_10__22_ ,
  \xz.mem_with_zero_10__21_ ,\xz.mem_with_zero_10__20_ ,\xz.mem_with_zero_10__19_ ,
  \xz.mem_with_zero_10__18_ ,\xz.mem_with_zero_10__17_ ,\xz.mem_with_zero_10__16_ ,
  \xz.mem_with_zero_10__15_ ,\xz.mem_with_zero_10__14_ ,\xz.mem_with_zero_10__13_ ,
  \xz.mem_with_zero_10__12_ ,\xz.mem_with_zero_10__11_ ,\xz.mem_with_zero_10__10_ ,
  \xz.mem_with_zero_10__9_ ,\xz.mem_with_zero_10__8_ ,\xz.mem_with_zero_10__7_ ,
  \xz.mem_with_zero_10__6_ ,\xz.mem_with_zero_10__5_ ,\xz.mem_with_zero_10__4_ ,
  \xz.mem_with_zero_10__3_ ,\xz.mem_with_zero_10__2_ ,\xz.mem_with_zero_10__1_ ,
  \xz.mem_with_zero_10__0_ ,\xz.mem_with_zero_9__31_ ,\xz.mem_with_zero_9__30_ ,
  \xz.mem_with_zero_9__29_ ,\xz.mem_with_zero_9__28_ ,\xz.mem_with_zero_9__27_ ,
  \xz.mem_with_zero_9__26_ ,\xz.mem_with_zero_9__25_ ,\xz.mem_with_zero_9__24_ ,
  \xz.mem_with_zero_9__23_ ,\xz.mem_with_zero_9__22_ ,\xz.mem_with_zero_9__21_ ,
  \xz.mem_with_zero_9__20_ ,\xz.mem_with_zero_9__19_ ,\xz.mem_with_zero_9__18_ ,
  \xz.mem_with_zero_9__17_ ,\xz.mem_with_zero_9__16_ ,\xz.mem_with_zero_9__15_ ,
  \xz.mem_with_zero_9__14_ ,\xz.mem_with_zero_9__13_ ,\xz.mem_with_zero_9__12_ ,
  \xz.mem_with_zero_9__11_ ,\xz.mem_with_zero_9__10_ ,\xz.mem_with_zero_9__9_ ,\xz.mem_with_zero_9__8_ ,
  \xz.mem_with_zero_9__7_ ,\xz.mem_with_zero_9__6_ ,\xz.mem_with_zero_9__5_ ,
  \xz.mem_with_zero_9__4_ ,\xz.mem_with_zero_9__3_ ,\xz.mem_with_zero_9__2_ ,
  \xz.mem_with_zero_9__1_ ,\xz.mem_with_zero_9__0_ ,\xz.mem_with_zero_8__31_ ,
  \xz.mem_with_zero_8__30_ ,\xz.mem_with_zero_8__29_ ,\xz.mem_with_zero_8__28_ ,
  \xz.mem_with_zero_8__27_ ,\xz.mem_with_zero_8__26_ ,\xz.mem_with_zero_8__25_ ,
  \xz.mem_with_zero_8__24_ ,\xz.mem_with_zero_8__23_ ,\xz.mem_with_zero_8__22_ ,
  \xz.mem_with_zero_8__21_ ,\xz.mem_with_zero_8__20_ ,\xz.mem_with_zero_8__19_ ,
  \xz.mem_with_zero_8__18_ ,\xz.mem_with_zero_8__17_ ,\xz.mem_with_zero_8__16_ ,\xz.mem_with_zero_8__15_ ,
  \xz.mem_with_zero_8__14_ ,\xz.mem_with_zero_8__13_ ,\xz.mem_with_zero_8__12_ ,
  \xz.mem_with_zero_8__11_ ,\xz.mem_with_zero_8__10_ ,\xz.mem_with_zero_8__9_ ,
  \xz.mem_with_zero_8__8_ ,\xz.mem_with_zero_8__7_ ,\xz.mem_with_zero_8__6_ ,
  \xz.mem_with_zero_8__5_ ,\xz.mem_with_zero_8__4_ ,\xz.mem_with_zero_8__3_ ,
  \xz.mem_with_zero_8__2_ ,\xz.mem_with_zero_8__1_ ,\xz.mem_with_zero_8__0_ ,
  \xz.mem_with_zero_7__31_ ,\xz.mem_with_zero_7__30_ ,\xz.mem_with_zero_7__29_ ,
  \xz.mem_with_zero_7__28_ ,\xz.mem_with_zero_7__27_ ,\xz.mem_with_zero_7__26_ ,
  \xz.mem_with_zero_7__25_ ,\xz.mem_with_zero_7__24_ ,\xz.mem_with_zero_7__23_ ,\xz.mem_with_zero_7__22_ ,
  \xz.mem_with_zero_7__21_ ,\xz.mem_with_zero_7__20_ ,\xz.mem_with_zero_7__19_ ,
  \xz.mem_with_zero_7__18_ ,\xz.mem_with_zero_7__17_ ,\xz.mem_with_zero_7__16_ ,
  \xz.mem_with_zero_7__15_ ,\xz.mem_with_zero_7__14_ ,\xz.mem_with_zero_7__13_ ,
  \xz.mem_with_zero_7__12_ ,\xz.mem_with_zero_7__11_ ,\xz.mem_with_zero_7__10_ ,
  \xz.mem_with_zero_7__9_ ,\xz.mem_with_zero_7__8_ ,\xz.mem_with_zero_7__7_ ,
  \xz.mem_with_zero_7__6_ ,\xz.mem_with_zero_7__5_ ,\xz.mem_with_zero_7__4_ ,
  \xz.mem_with_zero_7__3_ ,\xz.mem_with_zero_7__2_ ,\xz.mem_with_zero_7__1_ ,
  \xz.mem_with_zero_7__0_ ,\xz.mem_with_zero_6__31_ ,\xz.mem_with_zero_6__30_ ,\xz.mem_with_zero_6__29_ ,
  \xz.mem_with_zero_6__28_ ,\xz.mem_with_zero_6__27_ ,\xz.mem_with_zero_6__26_ ,
  \xz.mem_with_zero_6__25_ ,\xz.mem_with_zero_6__24_ ,\xz.mem_with_zero_6__23_ ,
  \xz.mem_with_zero_6__22_ ,\xz.mem_with_zero_6__21_ ,\xz.mem_with_zero_6__20_ ,
  \xz.mem_with_zero_6__19_ ,\xz.mem_with_zero_6__18_ ,\xz.mem_with_zero_6__17_ ,
  \xz.mem_with_zero_6__16_ ,\xz.mem_with_zero_6__15_ ,\xz.mem_with_zero_6__14_ ,
  \xz.mem_with_zero_6__13_ ,\xz.mem_with_zero_6__12_ ,\xz.mem_with_zero_6__11_ ,
  \xz.mem_with_zero_6__10_ ,\xz.mem_with_zero_6__9_ ,\xz.mem_with_zero_6__8_ ,
  \xz.mem_with_zero_6__7_ ,\xz.mem_with_zero_6__6_ ,\xz.mem_with_zero_6__5_ ,
  \xz.mem_with_zero_6__4_ ,\xz.mem_with_zero_6__3_ ,\xz.mem_with_zero_6__2_ ,\xz.mem_with_zero_6__1_ ,
  \xz.mem_with_zero_6__0_ ,\xz.mem_with_zero_5__31_ ,\xz.mem_with_zero_5__30_ ,
  \xz.mem_with_zero_5__29_ ,\xz.mem_with_zero_5__28_ ,\xz.mem_with_zero_5__27_ ,
  \xz.mem_with_zero_5__26_ ,\xz.mem_with_zero_5__25_ ,\xz.mem_with_zero_5__24_ ,
  \xz.mem_with_zero_5__23_ ,\xz.mem_with_zero_5__22_ ,\xz.mem_with_zero_5__21_ ,
  \xz.mem_with_zero_5__20_ ,\xz.mem_with_zero_5__19_ ,\xz.mem_with_zero_5__18_ ,
  \xz.mem_with_zero_5__17_ ,\xz.mem_with_zero_5__16_ ,\xz.mem_with_zero_5__15_ ,
  \xz.mem_with_zero_5__14_ ,\xz.mem_with_zero_5__13_ ,\xz.mem_with_zero_5__12_ ,
  \xz.mem_with_zero_5__11_ ,\xz.mem_with_zero_5__10_ ,\xz.mem_with_zero_5__9_ ,
  \xz.mem_with_zero_5__8_ ,\xz.mem_with_zero_5__7_ ,\xz.mem_with_zero_5__6_ ,\xz.mem_with_zero_5__5_ ,
  \xz.mem_with_zero_5__4_ ,\xz.mem_with_zero_5__3_ ,\xz.mem_with_zero_5__2_ ,
  \xz.mem_with_zero_5__1_ ,\xz.mem_with_zero_5__0_ ,\xz.mem_with_zero_4__31_ ,
  \xz.mem_with_zero_4__30_ ,\xz.mem_with_zero_4__29_ ,\xz.mem_with_zero_4__28_ ,
  \xz.mem_with_zero_4__27_ ,\xz.mem_with_zero_4__26_ ,\xz.mem_with_zero_4__25_ ,
  \xz.mem_with_zero_4__24_ ,\xz.mem_with_zero_4__23_ ,\xz.mem_with_zero_4__22_ ,
  \xz.mem_with_zero_4__21_ ,\xz.mem_with_zero_4__20_ ,\xz.mem_with_zero_4__19_ ,
  \xz.mem_with_zero_4__18_ ,\xz.mem_with_zero_4__17_ ,\xz.mem_with_zero_4__16_ ,
  \xz.mem_with_zero_4__15_ ,\xz.mem_with_zero_4__14_ ,\xz.mem_with_zero_4__13_ ,
  \xz.mem_with_zero_4__12_ ,\xz.mem_with_zero_4__11_ ,\xz.mem_with_zero_4__10_ ,
  \xz.mem_with_zero_4__9_ ,\xz.mem_with_zero_4__8_ ,\xz.mem_with_zero_4__7_ ,\xz.mem_with_zero_4__6_ ,
  \xz.mem_with_zero_4__5_ ,\xz.mem_with_zero_4__4_ ,\xz.mem_with_zero_4__3_ ,
  \xz.mem_with_zero_4__2_ ,\xz.mem_with_zero_4__1_ ,\xz.mem_with_zero_4__0_ ,
  \xz.mem_with_zero_3__31_ ,\xz.mem_with_zero_3__30_ ,\xz.mem_with_zero_3__29_ ,
  \xz.mem_with_zero_3__28_ ,\xz.mem_with_zero_3__27_ ,\xz.mem_with_zero_3__26_ ,
  \xz.mem_with_zero_3__25_ ,\xz.mem_with_zero_3__24_ ,\xz.mem_with_zero_3__23_ ,
  \xz.mem_with_zero_3__22_ ,\xz.mem_with_zero_3__21_ ,\xz.mem_with_zero_3__20_ ,
  \xz.mem_with_zero_3__19_ ,\xz.mem_with_zero_3__18_ ,\xz.mem_with_zero_3__17_ ,
  \xz.mem_with_zero_3__16_ ,\xz.mem_with_zero_3__15_ ,\xz.mem_with_zero_3__14_ ,
  \xz.mem_with_zero_3__13_ ,\xz.mem_with_zero_3__12_ ,\xz.mem_with_zero_3__11_ ,\xz.mem_with_zero_3__10_ ,
  \xz.mem_with_zero_3__9_ ,\xz.mem_with_zero_3__8_ ,\xz.mem_with_zero_3__7_ ,
  \xz.mem_with_zero_3__6_ ,\xz.mem_with_zero_3__5_ ,\xz.mem_with_zero_3__4_ ,
  \xz.mem_with_zero_3__3_ ,\xz.mem_with_zero_3__2_ ,\xz.mem_with_zero_3__1_ ,
  \xz.mem_with_zero_3__0_ ,\xz.mem_with_zero_2__31_ ,\xz.mem_with_zero_2__30_ ,
  \xz.mem_with_zero_2__29_ ,\xz.mem_with_zero_2__28_ ,\xz.mem_with_zero_2__27_ ,
  \xz.mem_with_zero_2__26_ ,\xz.mem_with_zero_2__25_ ,\xz.mem_with_zero_2__24_ ,
  \xz.mem_with_zero_2__23_ ,\xz.mem_with_zero_2__22_ ,\xz.mem_with_zero_2__21_ ,
  \xz.mem_with_zero_2__20_ ,\xz.mem_with_zero_2__19_ ,\xz.mem_with_zero_2__18_ ,\xz.mem_with_zero_2__17_ ,
  \xz.mem_with_zero_2__16_ ,\xz.mem_with_zero_2__15_ ,\xz.mem_with_zero_2__14_ ,
  \xz.mem_with_zero_2__13_ ,\xz.mem_with_zero_2__12_ ,\xz.mem_with_zero_2__11_ ,
  \xz.mem_with_zero_2__10_ ,\xz.mem_with_zero_2__9_ ,\xz.mem_with_zero_2__8_ ,
  \xz.mem_with_zero_2__7_ ,\xz.mem_with_zero_2__6_ ,\xz.mem_with_zero_2__5_ ,
  \xz.mem_with_zero_2__4_ ,\xz.mem_with_zero_2__3_ ,\xz.mem_with_zero_2__2_ ,
  \xz.mem_with_zero_2__1_ ,\xz.mem_with_zero_2__0_ ,\xz.mem_with_zero_1__31_ ,
  \xz.mem_with_zero_1__30_ ,\xz.mem_with_zero_1__29_ ,\xz.mem_with_zero_1__28_ ,
  \xz.mem_with_zero_1__27_ ,\xz.mem_with_zero_1__26_ ,\xz.mem_with_zero_1__25_ ,\xz.mem_with_zero_1__24_ ,
  \xz.mem_with_zero_1__23_ ,\xz.mem_with_zero_1__22_ ,\xz.mem_with_zero_1__21_ ,
  \xz.mem_with_zero_1__20_ ,\xz.mem_with_zero_1__19_ ,\xz.mem_with_zero_1__18_ ,
  \xz.mem_with_zero_1__17_ ,\xz.mem_with_zero_1__16_ ,\xz.mem_with_zero_1__15_ ,
  \xz.mem_with_zero_1__14_ ,\xz.mem_with_zero_1__13_ ,\xz.mem_with_zero_1__12_ ,
  \xz.mem_with_zero_1__11_ ,\xz.mem_with_zero_1__10_ ,\xz.mem_with_zero_1__9_ ,
  \xz.mem_with_zero_1__8_ ,\xz.mem_with_zero_1__7_ ,\xz.mem_with_zero_1__6_ ,
  \xz.mem_with_zero_1__5_ ,\xz.mem_with_zero_1__4_ ,\xz.mem_with_zero_1__3_ ,
  \xz.mem_with_zero_1__2_ ,\xz.mem_with_zero_1__1_ ,\xz.mem_with_zero_1__0_ ,N9,N10,N11,N12,N13,N14,N15,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,
  N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223;
  wire [9:0] r_addr_r;
  reg r_addr_r_9_sv2v_reg,r_addr_r_8_sv2v_reg,r_addr_r_7_sv2v_reg,r_addr_r_6_sv2v_reg,
  r_addr_r_5_sv2v_reg,r_addr_r_4_sv2v_reg,r_addr_r_3_sv2v_reg,r_addr_r_2_sv2v_reg,
  r_addr_r_1_sv2v_reg,r_addr_r_0_sv2v_reg,\xz.mem_with_zero_31__31__sv2v_reg ,
  \xz.mem_with_zero_31__30__sv2v_reg ,\xz.mem_with_zero_31__29__sv2v_reg ,
  \xz.mem_with_zero_31__28__sv2v_reg ,\xz.mem_with_zero_31__27__sv2v_reg ,
  \xz.mem_with_zero_31__26__sv2v_reg ,\xz.mem_with_zero_31__25__sv2v_reg ,
  \xz.mem_with_zero_31__24__sv2v_reg ,\xz.mem_with_zero_31__23__sv2v_reg ,\xz.mem_with_zero_31__22__sv2v_reg ,
  \xz.mem_with_zero_31__21__sv2v_reg ,\xz.mem_with_zero_31__20__sv2v_reg ,
  \xz.mem_with_zero_31__19__sv2v_reg ,\xz.mem_with_zero_31__18__sv2v_reg ,
  \xz.mem_with_zero_31__17__sv2v_reg ,\xz.mem_with_zero_31__16__sv2v_reg ,
  \xz.mem_with_zero_31__15__sv2v_reg ,\xz.mem_with_zero_31__14__sv2v_reg ,
  \xz.mem_with_zero_31__13__sv2v_reg ,\xz.mem_with_zero_31__12__sv2v_reg ,\xz.mem_with_zero_31__11__sv2v_reg ,
  \xz.mem_with_zero_31__10__sv2v_reg ,\xz.mem_with_zero_31__9__sv2v_reg ,
  \xz.mem_with_zero_31__8__sv2v_reg ,\xz.mem_with_zero_31__7__sv2v_reg ,
  \xz.mem_with_zero_31__6__sv2v_reg ,\xz.mem_with_zero_31__5__sv2v_reg ,
  \xz.mem_with_zero_31__4__sv2v_reg ,\xz.mem_with_zero_31__3__sv2v_reg ,\xz.mem_with_zero_31__2__sv2v_reg ,
  \xz.mem_with_zero_31__1__sv2v_reg ,\xz.mem_with_zero_31__0__sv2v_reg ,
  \xz.mem_with_zero_30__31__sv2v_reg ,\xz.mem_with_zero_30__30__sv2v_reg ,
  \xz.mem_with_zero_30__29__sv2v_reg ,\xz.mem_with_zero_30__28__sv2v_reg ,
  \xz.mem_with_zero_30__27__sv2v_reg ,\xz.mem_with_zero_30__26__sv2v_reg ,\xz.mem_with_zero_30__25__sv2v_reg ,
  \xz.mem_with_zero_30__24__sv2v_reg ,\xz.mem_with_zero_30__23__sv2v_reg ,
  \xz.mem_with_zero_30__22__sv2v_reg ,\xz.mem_with_zero_30__21__sv2v_reg ,
  \xz.mem_with_zero_30__20__sv2v_reg ,\xz.mem_with_zero_30__19__sv2v_reg ,
  \xz.mem_with_zero_30__18__sv2v_reg ,\xz.mem_with_zero_30__17__sv2v_reg ,\xz.mem_with_zero_30__16__sv2v_reg ,
  \xz.mem_with_zero_30__15__sv2v_reg ,\xz.mem_with_zero_30__14__sv2v_reg ,
  \xz.mem_with_zero_30__13__sv2v_reg ,\xz.mem_with_zero_30__12__sv2v_reg ,
  \xz.mem_with_zero_30__11__sv2v_reg ,\xz.mem_with_zero_30__10__sv2v_reg ,
  \xz.mem_with_zero_30__9__sv2v_reg ,\xz.mem_with_zero_30__8__sv2v_reg ,\xz.mem_with_zero_30__7__sv2v_reg ,
  \xz.mem_with_zero_30__6__sv2v_reg ,\xz.mem_with_zero_30__5__sv2v_reg ,
  \xz.mem_with_zero_30__4__sv2v_reg ,\xz.mem_with_zero_30__3__sv2v_reg ,
  \xz.mem_with_zero_30__2__sv2v_reg ,\xz.mem_with_zero_30__1__sv2v_reg ,
  \xz.mem_with_zero_30__0__sv2v_reg ,\xz.mem_with_zero_29__31__sv2v_reg ,\xz.mem_with_zero_29__30__sv2v_reg ,
  \xz.mem_with_zero_29__29__sv2v_reg ,\xz.mem_with_zero_29__28__sv2v_reg ,
  \xz.mem_with_zero_29__27__sv2v_reg ,\xz.mem_with_zero_29__26__sv2v_reg ,
  \xz.mem_with_zero_29__25__sv2v_reg ,\xz.mem_with_zero_29__24__sv2v_reg ,
  \xz.mem_with_zero_29__23__sv2v_reg ,\xz.mem_with_zero_29__22__sv2v_reg ,\xz.mem_with_zero_29__21__sv2v_reg ,
  \xz.mem_with_zero_29__20__sv2v_reg ,\xz.mem_with_zero_29__19__sv2v_reg ,
  \xz.mem_with_zero_29__18__sv2v_reg ,\xz.mem_with_zero_29__17__sv2v_reg ,
  \xz.mem_with_zero_29__16__sv2v_reg ,\xz.mem_with_zero_29__15__sv2v_reg ,
  \xz.mem_with_zero_29__14__sv2v_reg ,\xz.mem_with_zero_29__13__sv2v_reg ,
  \xz.mem_with_zero_29__12__sv2v_reg ,\xz.mem_with_zero_29__11__sv2v_reg ,\xz.mem_with_zero_29__10__sv2v_reg ,
  \xz.mem_with_zero_29__9__sv2v_reg ,\xz.mem_with_zero_29__8__sv2v_reg ,
  \xz.mem_with_zero_29__7__sv2v_reg ,\xz.mem_with_zero_29__6__sv2v_reg ,
  \xz.mem_with_zero_29__5__sv2v_reg ,\xz.mem_with_zero_29__4__sv2v_reg ,
  \xz.mem_with_zero_29__3__sv2v_reg ,\xz.mem_with_zero_29__2__sv2v_reg ,\xz.mem_with_zero_29__1__sv2v_reg ,
  \xz.mem_with_zero_29__0__sv2v_reg ,\xz.mem_with_zero_28__31__sv2v_reg ,
  \xz.mem_with_zero_28__30__sv2v_reg ,\xz.mem_with_zero_28__29__sv2v_reg ,
  \xz.mem_with_zero_28__28__sv2v_reg ,\xz.mem_with_zero_28__27__sv2v_reg ,
  \xz.mem_with_zero_28__26__sv2v_reg ,\xz.mem_with_zero_28__25__sv2v_reg ,\xz.mem_with_zero_28__24__sv2v_reg ,
  \xz.mem_with_zero_28__23__sv2v_reg ,\xz.mem_with_zero_28__22__sv2v_reg ,
  \xz.mem_with_zero_28__21__sv2v_reg ,\xz.mem_with_zero_28__20__sv2v_reg ,
  \xz.mem_with_zero_28__19__sv2v_reg ,\xz.mem_with_zero_28__18__sv2v_reg ,
  \xz.mem_with_zero_28__17__sv2v_reg ,\xz.mem_with_zero_28__16__sv2v_reg ,\xz.mem_with_zero_28__15__sv2v_reg ,
  \xz.mem_with_zero_28__14__sv2v_reg ,\xz.mem_with_zero_28__13__sv2v_reg ,
  \xz.mem_with_zero_28__12__sv2v_reg ,\xz.mem_with_zero_28__11__sv2v_reg ,
  \xz.mem_with_zero_28__10__sv2v_reg ,\xz.mem_with_zero_28__9__sv2v_reg ,
  \xz.mem_with_zero_28__8__sv2v_reg ,\xz.mem_with_zero_28__7__sv2v_reg ,\xz.mem_with_zero_28__6__sv2v_reg ,
  \xz.mem_with_zero_28__5__sv2v_reg ,\xz.mem_with_zero_28__4__sv2v_reg ,
  \xz.mem_with_zero_28__3__sv2v_reg ,\xz.mem_with_zero_28__2__sv2v_reg ,
  \xz.mem_with_zero_28__1__sv2v_reg ,\xz.mem_with_zero_28__0__sv2v_reg ,
  \xz.mem_with_zero_27__31__sv2v_reg ,\xz.mem_with_zero_27__30__sv2v_reg ,\xz.mem_with_zero_27__29__sv2v_reg ,
  \xz.mem_with_zero_27__28__sv2v_reg ,\xz.mem_with_zero_27__27__sv2v_reg ,
  \xz.mem_with_zero_27__26__sv2v_reg ,\xz.mem_with_zero_27__25__sv2v_reg ,
  \xz.mem_with_zero_27__24__sv2v_reg ,\xz.mem_with_zero_27__23__sv2v_reg ,
  \xz.mem_with_zero_27__22__sv2v_reg ,\xz.mem_with_zero_27__21__sv2v_reg ,\xz.mem_with_zero_27__20__sv2v_reg ,
  \xz.mem_with_zero_27__19__sv2v_reg ,\xz.mem_with_zero_27__18__sv2v_reg ,
  \xz.mem_with_zero_27__17__sv2v_reg ,\xz.mem_with_zero_27__16__sv2v_reg ,
  \xz.mem_with_zero_27__15__sv2v_reg ,\xz.mem_with_zero_27__14__sv2v_reg ,
  \xz.mem_with_zero_27__13__sv2v_reg ,\xz.mem_with_zero_27__12__sv2v_reg ,
  \xz.mem_with_zero_27__11__sv2v_reg ,\xz.mem_with_zero_27__10__sv2v_reg ,\xz.mem_with_zero_27__9__sv2v_reg ,
  \xz.mem_with_zero_27__8__sv2v_reg ,\xz.mem_with_zero_27__7__sv2v_reg ,
  \xz.mem_with_zero_27__6__sv2v_reg ,\xz.mem_with_zero_27__5__sv2v_reg ,
  \xz.mem_with_zero_27__4__sv2v_reg ,\xz.mem_with_zero_27__3__sv2v_reg ,\xz.mem_with_zero_27__2__sv2v_reg ,
  \xz.mem_with_zero_27__1__sv2v_reg ,\xz.mem_with_zero_27__0__sv2v_reg ,
  \xz.mem_with_zero_26__31__sv2v_reg ,\xz.mem_with_zero_26__30__sv2v_reg ,
  \xz.mem_with_zero_26__29__sv2v_reg ,\xz.mem_with_zero_26__28__sv2v_reg ,
  \xz.mem_with_zero_26__27__sv2v_reg ,\xz.mem_with_zero_26__26__sv2v_reg ,
  \xz.mem_with_zero_26__25__sv2v_reg ,\xz.mem_with_zero_26__24__sv2v_reg ,\xz.mem_with_zero_26__23__sv2v_reg ,
  \xz.mem_with_zero_26__22__sv2v_reg ,\xz.mem_with_zero_26__21__sv2v_reg ,
  \xz.mem_with_zero_26__20__sv2v_reg ,\xz.mem_with_zero_26__19__sv2v_reg ,
  \xz.mem_with_zero_26__18__sv2v_reg ,\xz.mem_with_zero_26__17__sv2v_reg ,
  \xz.mem_with_zero_26__16__sv2v_reg ,\xz.mem_with_zero_26__15__sv2v_reg ,\xz.mem_with_zero_26__14__sv2v_reg ,
  \xz.mem_with_zero_26__13__sv2v_reg ,\xz.mem_with_zero_26__12__sv2v_reg ,
  \xz.mem_with_zero_26__11__sv2v_reg ,\xz.mem_with_zero_26__10__sv2v_reg ,
  \xz.mem_with_zero_26__9__sv2v_reg ,\xz.mem_with_zero_26__8__sv2v_reg ,
  \xz.mem_with_zero_26__7__sv2v_reg ,\xz.mem_with_zero_26__6__sv2v_reg ,\xz.mem_with_zero_26__5__sv2v_reg ,
  \xz.mem_with_zero_26__4__sv2v_reg ,\xz.mem_with_zero_26__3__sv2v_reg ,
  \xz.mem_with_zero_26__2__sv2v_reg ,\xz.mem_with_zero_26__1__sv2v_reg ,
  \xz.mem_with_zero_26__0__sv2v_reg ,\xz.mem_with_zero_25__31__sv2v_reg ,
  \xz.mem_with_zero_25__30__sv2v_reg ,\xz.mem_with_zero_25__29__sv2v_reg ,\xz.mem_with_zero_25__28__sv2v_reg ,
  \xz.mem_with_zero_25__27__sv2v_reg ,\xz.mem_with_zero_25__26__sv2v_reg ,
  \xz.mem_with_zero_25__25__sv2v_reg ,\xz.mem_with_zero_25__24__sv2v_reg ,
  \xz.mem_with_zero_25__23__sv2v_reg ,\xz.mem_with_zero_25__22__sv2v_reg ,
  \xz.mem_with_zero_25__21__sv2v_reg ,\xz.mem_with_zero_25__20__sv2v_reg ,\xz.mem_with_zero_25__19__sv2v_reg ,
  \xz.mem_with_zero_25__18__sv2v_reg ,\xz.mem_with_zero_25__17__sv2v_reg ,
  \xz.mem_with_zero_25__16__sv2v_reg ,\xz.mem_with_zero_25__15__sv2v_reg ,
  \xz.mem_with_zero_25__14__sv2v_reg ,\xz.mem_with_zero_25__13__sv2v_reg ,
  \xz.mem_with_zero_25__12__sv2v_reg ,\xz.mem_with_zero_25__11__sv2v_reg ,
  \xz.mem_with_zero_25__10__sv2v_reg ,\xz.mem_with_zero_25__9__sv2v_reg ,\xz.mem_with_zero_25__8__sv2v_reg ,
  \xz.mem_with_zero_25__7__sv2v_reg ,\xz.mem_with_zero_25__6__sv2v_reg ,
  \xz.mem_with_zero_25__5__sv2v_reg ,\xz.mem_with_zero_25__4__sv2v_reg ,
  \xz.mem_with_zero_25__3__sv2v_reg ,\xz.mem_with_zero_25__2__sv2v_reg ,\xz.mem_with_zero_25__1__sv2v_reg ,
  \xz.mem_with_zero_25__0__sv2v_reg ,\xz.mem_with_zero_24__31__sv2v_reg ,
  \xz.mem_with_zero_24__30__sv2v_reg ,\xz.mem_with_zero_24__29__sv2v_reg ,
  \xz.mem_with_zero_24__28__sv2v_reg ,\xz.mem_with_zero_24__27__sv2v_reg ,
  \xz.mem_with_zero_24__26__sv2v_reg ,\xz.mem_with_zero_24__25__sv2v_reg ,
  \xz.mem_with_zero_24__24__sv2v_reg ,\xz.mem_with_zero_24__23__sv2v_reg ,\xz.mem_with_zero_24__22__sv2v_reg ,
  \xz.mem_with_zero_24__21__sv2v_reg ,\xz.mem_with_zero_24__20__sv2v_reg ,
  \xz.mem_with_zero_24__19__sv2v_reg ,\xz.mem_with_zero_24__18__sv2v_reg ,
  \xz.mem_with_zero_24__17__sv2v_reg ,\xz.mem_with_zero_24__16__sv2v_reg ,
  \xz.mem_with_zero_24__15__sv2v_reg ,\xz.mem_with_zero_24__14__sv2v_reg ,\xz.mem_with_zero_24__13__sv2v_reg ,
  \xz.mem_with_zero_24__12__sv2v_reg ,\xz.mem_with_zero_24__11__sv2v_reg ,
  \xz.mem_with_zero_24__10__sv2v_reg ,\xz.mem_with_zero_24__9__sv2v_reg ,
  \xz.mem_with_zero_24__8__sv2v_reg ,\xz.mem_with_zero_24__7__sv2v_reg ,
  \xz.mem_with_zero_24__6__sv2v_reg ,\xz.mem_with_zero_24__5__sv2v_reg ,\xz.mem_with_zero_24__4__sv2v_reg ,
  \xz.mem_with_zero_24__3__sv2v_reg ,\xz.mem_with_zero_24__2__sv2v_reg ,
  \xz.mem_with_zero_24__1__sv2v_reg ,\xz.mem_with_zero_24__0__sv2v_reg ,
  \xz.mem_with_zero_23__31__sv2v_reg ,\xz.mem_with_zero_23__30__sv2v_reg ,
  \xz.mem_with_zero_23__29__sv2v_reg ,\xz.mem_with_zero_23__28__sv2v_reg ,\xz.mem_with_zero_23__27__sv2v_reg ,
  \xz.mem_with_zero_23__26__sv2v_reg ,\xz.mem_with_zero_23__25__sv2v_reg ,
  \xz.mem_with_zero_23__24__sv2v_reg ,\xz.mem_with_zero_23__23__sv2v_reg ,
  \xz.mem_with_zero_23__22__sv2v_reg ,\xz.mem_with_zero_23__21__sv2v_reg ,
  \xz.mem_with_zero_23__20__sv2v_reg ,\xz.mem_with_zero_23__19__sv2v_reg ,\xz.mem_with_zero_23__18__sv2v_reg ,
  \xz.mem_with_zero_23__17__sv2v_reg ,\xz.mem_with_zero_23__16__sv2v_reg ,
  \xz.mem_with_zero_23__15__sv2v_reg ,\xz.mem_with_zero_23__14__sv2v_reg ,
  \xz.mem_with_zero_23__13__sv2v_reg ,\xz.mem_with_zero_23__12__sv2v_reg ,
  \xz.mem_with_zero_23__11__sv2v_reg ,\xz.mem_with_zero_23__10__sv2v_reg ,
  \xz.mem_with_zero_23__9__sv2v_reg ,\xz.mem_with_zero_23__8__sv2v_reg ,\xz.mem_with_zero_23__7__sv2v_reg ,
  \xz.mem_with_zero_23__6__sv2v_reg ,\xz.mem_with_zero_23__5__sv2v_reg ,
  \xz.mem_with_zero_23__4__sv2v_reg ,\xz.mem_with_zero_23__3__sv2v_reg ,
  \xz.mem_with_zero_23__2__sv2v_reg ,\xz.mem_with_zero_23__1__sv2v_reg ,\xz.mem_with_zero_23__0__sv2v_reg ,
  \xz.mem_with_zero_22__31__sv2v_reg ,\xz.mem_with_zero_22__30__sv2v_reg ,
  \xz.mem_with_zero_22__29__sv2v_reg ,\xz.mem_with_zero_22__28__sv2v_reg ,
  \xz.mem_with_zero_22__27__sv2v_reg ,\xz.mem_with_zero_22__26__sv2v_reg ,
  \xz.mem_with_zero_22__25__sv2v_reg ,\xz.mem_with_zero_22__24__sv2v_reg ,
  \xz.mem_with_zero_22__23__sv2v_reg ,\xz.mem_with_zero_22__22__sv2v_reg ,\xz.mem_with_zero_22__21__sv2v_reg ,
  \xz.mem_with_zero_22__20__sv2v_reg ,\xz.mem_with_zero_22__19__sv2v_reg ,
  \xz.mem_with_zero_22__18__sv2v_reg ,\xz.mem_with_zero_22__17__sv2v_reg ,
  \xz.mem_with_zero_22__16__sv2v_reg ,\xz.mem_with_zero_22__15__sv2v_reg ,
  \xz.mem_with_zero_22__14__sv2v_reg ,\xz.mem_with_zero_22__13__sv2v_reg ,\xz.mem_with_zero_22__12__sv2v_reg ,
  \xz.mem_with_zero_22__11__sv2v_reg ,\xz.mem_with_zero_22__10__sv2v_reg ,
  \xz.mem_with_zero_22__9__sv2v_reg ,\xz.mem_with_zero_22__8__sv2v_reg ,
  \xz.mem_with_zero_22__7__sv2v_reg ,\xz.mem_with_zero_22__6__sv2v_reg ,
  \xz.mem_with_zero_22__5__sv2v_reg ,\xz.mem_with_zero_22__4__sv2v_reg ,\xz.mem_with_zero_22__3__sv2v_reg ,
  \xz.mem_with_zero_22__2__sv2v_reg ,\xz.mem_with_zero_22__1__sv2v_reg ,
  \xz.mem_with_zero_22__0__sv2v_reg ,\xz.mem_with_zero_21__31__sv2v_reg ,
  \xz.mem_with_zero_21__30__sv2v_reg ,\xz.mem_with_zero_21__29__sv2v_reg ,
  \xz.mem_with_zero_21__28__sv2v_reg ,\xz.mem_with_zero_21__27__sv2v_reg ,\xz.mem_with_zero_21__26__sv2v_reg ,
  \xz.mem_with_zero_21__25__sv2v_reg ,\xz.mem_with_zero_21__24__sv2v_reg ,
  \xz.mem_with_zero_21__23__sv2v_reg ,\xz.mem_with_zero_21__22__sv2v_reg ,
  \xz.mem_with_zero_21__21__sv2v_reg ,\xz.mem_with_zero_21__20__sv2v_reg ,
  \xz.mem_with_zero_21__19__sv2v_reg ,\xz.mem_with_zero_21__18__sv2v_reg ,\xz.mem_with_zero_21__17__sv2v_reg ,
  \xz.mem_with_zero_21__16__sv2v_reg ,\xz.mem_with_zero_21__15__sv2v_reg ,
  \xz.mem_with_zero_21__14__sv2v_reg ,\xz.mem_with_zero_21__13__sv2v_reg ,
  \xz.mem_with_zero_21__12__sv2v_reg ,\xz.mem_with_zero_21__11__sv2v_reg ,
  \xz.mem_with_zero_21__10__sv2v_reg ,\xz.mem_with_zero_21__9__sv2v_reg ,
  \xz.mem_with_zero_21__8__sv2v_reg ,\xz.mem_with_zero_21__7__sv2v_reg ,\xz.mem_with_zero_21__6__sv2v_reg ,
  \xz.mem_with_zero_21__5__sv2v_reg ,\xz.mem_with_zero_21__4__sv2v_reg ,
  \xz.mem_with_zero_21__3__sv2v_reg ,\xz.mem_with_zero_21__2__sv2v_reg ,
  \xz.mem_with_zero_21__1__sv2v_reg ,\xz.mem_with_zero_21__0__sv2v_reg ,\xz.mem_with_zero_20__31__sv2v_reg ,
  \xz.mem_with_zero_20__30__sv2v_reg ,\xz.mem_with_zero_20__29__sv2v_reg ,
  \xz.mem_with_zero_20__28__sv2v_reg ,\xz.mem_with_zero_20__27__sv2v_reg ,
  \xz.mem_with_zero_20__26__sv2v_reg ,\xz.mem_with_zero_20__25__sv2v_reg ,
  \xz.mem_with_zero_20__24__sv2v_reg ,\xz.mem_with_zero_20__23__sv2v_reg ,
  \xz.mem_with_zero_20__22__sv2v_reg ,\xz.mem_with_zero_20__21__sv2v_reg ,\xz.mem_with_zero_20__20__sv2v_reg ,
  \xz.mem_with_zero_20__19__sv2v_reg ,\xz.mem_with_zero_20__18__sv2v_reg ,
  \xz.mem_with_zero_20__17__sv2v_reg ,\xz.mem_with_zero_20__16__sv2v_reg ,
  \xz.mem_with_zero_20__15__sv2v_reg ,\xz.mem_with_zero_20__14__sv2v_reg ,
  \xz.mem_with_zero_20__13__sv2v_reg ,\xz.mem_with_zero_20__12__sv2v_reg ,\xz.mem_with_zero_20__11__sv2v_reg ,
  \xz.mem_with_zero_20__10__sv2v_reg ,\xz.mem_with_zero_20__9__sv2v_reg ,
  \xz.mem_with_zero_20__8__sv2v_reg ,\xz.mem_with_zero_20__7__sv2v_reg ,
  \xz.mem_with_zero_20__6__sv2v_reg ,\xz.mem_with_zero_20__5__sv2v_reg ,
  \xz.mem_with_zero_20__4__sv2v_reg ,\xz.mem_with_zero_20__3__sv2v_reg ,\xz.mem_with_zero_20__2__sv2v_reg ,
  \xz.mem_with_zero_20__1__sv2v_reg ,\xz.mem_with_zero_20__0__sv2v_reg ,
  \xz.mem_with_zero_19__31__sv2v_reg ,\xz.mem_with_zero_19__30__sv2v_reg ,
  \xz.mem_with_zero_19__29__sv2v_reg ,\xz.mem_with_zero_19__28__sv2v_reg ,
  \xz.mem_with_zero_19__27__sv2v_reg ,\xz.mem_with_zero_19__26__sv2v_reg ,\xz.mem_with_zero_19__25__sv2v_reg ,
  \xz.mem_with_zero_19__24__sv2v_reg ,\xz.mem_with_zero_19__23__sv2v_reg ,
  \xz.mem_with_zero_19__22__sv2v_reg ,\xz.mem_with_zero_19__21__sv2v_reg ,
  \xz.mem_with_zero_19__20__sv2v_reg ,\xz.mem_with_zero_19__19__sv2v_reg ,
  \xz.mem_with_zero_19__18__sv2v_reg ,\xz.mem_with_zero_19__17__sv2v_reg ,\xz.mem_with_zero_19__16__sv2v_reg ,
  \xz.mem_with_zero_19__15__sv2v_reg ,\xz.mem_with_zero_19__14__sv2v_reg ,
  \xz.mem_with_zero_19__13__sv2v_reg ,\xz.mem_with_zero_19__12__sv2v_reg ,
  \xz.mem_with_zero_19__11__sv2v_reg ,\xz.mem_with_zero_19__10__sv2v_reg ,
  \xz.mem_with_zero_19__9__sv2v_reg ,\xz.mem_with_zero_19__8__sv2v_reg ,
  \xz.mem_with_zero_19__7__sv2v_reg ,\xz.mem_with_zero_19__6__sv2v_reg ,\xz.mem_with_zero_19__5__sv2v_reg ,
  \xz.mem_with_zero_19__4__sv2v_reg ,\xz.mem_with_zero_19__3__sv2v_reg ,
  \xz.mem_with_zero_19__2__sv2v_reg ,\xz.mem_with_zero_19__1__sv2v_reg ,
  \xz.mem_with_zero_19__0__sv2v_reg ,\xz.mem_with_zero_18__31__sv2v_reg ,\xz.mem_with_zero_18__30__sv2v_reg ,
  \xz.mem_with_zero_18__29__sv2v_reg ,\xz.mem_with_zero_18__28__sv2v_reg ,
  \xz.mem_with_zero_18__27__sv2v_reg ,\xz.mem_with_zero_18__26__sv2v_reg ,
  \xz.mem_with_zero_18__25__sv2v_reg ,\xz.mem_with_zero_18__24__sv2v_reg ,
  \xz.mem_with_zero_18__23__sv2v_reg ,\xz.mem_with_zero_18__22__sv2v_reg ,
  \xz.mem_with_zero_18__21__sv2v_reg ,\xz.mem_with_zero_18__20__sv2v_reg ,\xz.mem_with_zero_18__19__sv2v_reg ,
  \xz.mem_with_zero_18__18__sv2v_reg ,\xz.mem_with_zero_18__17__sv2v_reg ,
  \xz.mem_with_zero_18__16__sv2v_reg ,\xz.mem_with_zero_18__15__sv2v_reg ,
  \xz.mem_with_zero_18__14__sv2v_reg ,\xz.mem_with_zero_18__13__sv2v_reg ,
  \xz.mem_with_zero_18__12__sv2v_reg ,\xz.mem_with_zero_18__11__sv2v_reg ,\xz.mem_with_zero_18__10__sv2v_reg ,
  \xz.mem_with_zero_18__9__sv2v_reg ,\xz.mem_with_zero_18__8__sv2v_reg ,
  \xz.mem_with_zero_18__7__sv2v_reg ,\xz.mem_with_zero_18__6__sv2v_reg ,
  \xz.mem_with_zero_18__5__sv2v_reg ,\xz.mem_with_zero_18__4__sv2v_reg ,
  \xz.mem_with_zero_18__3__sv2v_reg ,\xz.mem_with_zero_18__2__sv2v_reg ,\xz.mem_with_zero_18__1__sv2v_reg ,
  \xz.mem_with_zero_18__0__sv2v_reg ,\xz.mem_with_zero_17__31__sv2v_reg ,
  \xz.mem_with_zero_17__30__sv2v_reg ,\xz.mem_with_zero_17__29__sv2v_reg ,
  \xz.mem_with_zero_17__28__sv2v_reg ,\xz.mem_with_zero_17__27__sv2v_reg ,
  \xz.mem_with_zero_17__26__sv2v_reg ,\xz.mem_with_zero_17__25__sv2v_reg ,\xz.mem_with_zero_17__24__sv2v_reg ,
  \xz.mem_with_zero_17__23__sv2v_reg ,\xz.mem_with_zero_17__22__sv2v_reg ,
  \xz.mem_with_zero_17__21__sv2v_reg ,\xz.mem_with_zero_17__20__sv2v_reg ,
  \xz.mem_with_zero_17__19__sv2v_reg ,\xz.mem_with_zero_17__18__sv2v_reg ,
  \xz.mem_with_zero_17__17__sv2v_reg ,\xz.mem_with_zero_17__16__sv2v_reg ,\xz.mem_with_zero_17__15__sv2v_reg ,
  \xz.mem_with_zero_17__14__sv2v_reg ,\xz.mem_with_zero_17__13__sv2v_reg ,
  \xz.mem_with_zero_17__12__sv2v_reg ,\xz.mem_with_zero_17__11__sv2v_reg ,
  \xz.mem_with_zero_17__10__sv2v_reg ,\xz.mem_with_zero_17__9__sv2v_reg ,
  \xz.mem_with_zero_17__8__sv2v_reg ,\xz.mem_with_zero_17__7__sv2v_reg ,\xz.mem_with_zero_17__6__sv2v_reg ,
  \xz.mem_with_zero_17__5__sv2v_reg ,\xz.mem_with_zero_17__4__sv2v_reg ,
  \xz.mem_with_zero_17__3__sv2v_reg ,\xz.mem_with_zero_17__2__sv2v_reg ,
  \xz.mem_with_zero_17__1__sv2v_reg ,\xz.mem_with_zero_17__0__sv2v_reg ,
  \xz.mem_with_zero_16__31__sv2v_reg ,\xz.mem_with_zero_16__30__sv2v_reg ,\xz.mem_with_zero_16__29__sv2v_reg ,
  \xz.mem_with_zero_16__28__sv2v_reg ,\xz.mem_with_zero_16__27__sv2v_reg ,
  \xz.mem_with_zero_16__26__sv2v_reg ,\xz.mem_with_zero_16__25__sv2v_reg ,
  \xz.mem_with_zero_16__24__sv2v_reg ,\xz.mem_with_zero_16__23__sv2v_reg ,
  \xz.mem_with_zero_16__22__sv2v_reg ,\xz.mem_with_zero_16__21__sv2v_reg ,
  \xz.mem_with_zero_16__20__sv2v_reg ,\xz.mem_with_zero_16__19__sv2v_reg ,\xz.mem_with_zero_16__18__sv2v_reg ,
  \xz.mem_with_zero_16__17__sv2v_reg ,\xz.mem_with_zero_16__16__sv2v_reg ,
  \xz.mem_with_zero_16__15__sv2v_reg ,\xz.mem_with_zero_16__14__sv2v_reg ,
  \xz.mem_with_zero_16__13__sv2v_reg ,\xz.mem_with_zero_16__12__sv2v_reg ,
  \xz.mem_with_zero_16__11__sv2v_reg ,\xz.mem_with_zero_16__10__sv2v_reg ,\xz.mem_with_zero_16__9__sv2v_reg ,
  \xz.mem_with_zero_16__8__sv2v_reg ,\xz.mem_with_zero_16__7__sv2v_reg ,
  \xz.mem_with_zero_16__6__sv2v_reg ,\xz.mem_with_zero_16__5__sv2v_reg ,
  \xz.mem_with_zero_16__4__sv2v_reg ,\xz.mem_with_zero_16__3__sv2v_reg ,
  \xz.mem_with_zero_16__2__sv2v_reg ,\xz.mem_with_zero_16__1__sv2v_reg ,\xz.mem_with_zero_16__0__sv2v_reg ,
  \xz.mem_with_zero_15__31__sv2v_reg ,\xz.mem_with_zero_15__30__sv2v_reg ,
  \xz.mem_with_zero_15__29__sv2v_reg ,\xz.mem_with_zero_15__28__sv2v_reg ,
  \xz.mem_with_zero_15__27__sv2v_reg ,\xz.mem_with_zero_15__26__sv2v_reg ,
  \xz.mem_with_zero_15__25__sv2v_reg ,\xz.mem_with_zero_15__24__sv2v_reg ,\xz.mem_with_zero_15__23__sv2v_reg ,
  \xz.mem_with_zero_15__22__sv2v_reg ,\xz.mem_with_zero_15__21__sv2v_reg ,
  \xz.mem_with_zero_15__20__sv2v_reg ,\xz.mem_with_zero_15__19__sv2v_reg ,
  \xz.mem_with_zero_15__18__sv2v_reg ,\xz.mem_with_zero_15__17__sv2v_reg ,
  \xz.mem_with_zero_15__16__sv2v_reg ,\xz.mem_with_zero_15__15__sv2v_reg ,\xz.mem_with_zero_15__14__sv2v_reg ,
  \xz.mem_with_zero_15__13__sv2v_reg ,\xz.mem_with_zero_15__12__sv2v_reg ,
  \xz.mem_with_zero_15__11__sv2v_reg ,\xz.mem_with_zero_15__10__sv2v_reg ,
  \xz.mem_with_zero_15__9__sv2v_reg ,\xz.mem_with_zero_15__8__sv2v_reg ,
  \xz.mem_with_zero_15__7__sv2v_reg ,\xz.mem_with_zero_15__6__sv2v_reg ,\xz.mem_with_zero_15__5__sv2v_reg ,
  \xz.mem_with_zero_15__4__sv2v_reg ,\xz.mem_with_zero_15__3__sv2v_reg ,
  \xz.mem_with_zero_15__2__sv2v_reg ,\xz.mem_with_zero_15__1__sv2v_reg ,
  \xz.mem_with_zero_15__0__sv2v_reg ,\xz.mem_with_zero_14__31__sv2v_reg ,
  \xz.mem_with_zero_14__30__sv2v_reg ,\xz.mem_with_zero_14__29__sv2v_reg ,\xz.mem_with_zero_14__28__sv2v_reg ,
  \xz.mem_with_zero_14__27__sv2v_reg ,\xz.mem_with_zero_14__26__sv2v_reg ,
  \xz.mem_with_zero_14__25__sv2v_reg ,\xz.mem_with_zero_14__24__sv2v_reg ,
  \xz.mem_with_zero_14__23__sv2v_reg ,\xz.mem_with_zero_14__22__sv2v_reg ,
  \xz.mem_with_zero_14__21__sv2v_reg ,\xz.mem_with_zero_14__20__sv2v_reg ,
  \xz.mem_with_zero_14__19__sv2v_reg ,\xz.mem_with_zero_14__18__sv2v_reg ,\xz.mem_with_zero_14__17__sv2v_reg ,
  \xz.mem_with_zero_14__16__sv2v_reg ,\xz.mem_with_zero_14__15__sv2v_reg ,
  \xz.mem_with_zero_14__14__sv2v_reg ,\xz.mem_with_zero_14__13__sv2v_reg ,
  \xz.mem_with_zero_14__12__sv2v_reg ,\xz.mem_with_zero_14__11__sv2v_reg ,
  \xz.mem_with_zero_14__10__sv2v_reg ,\xz.mem_with_zero_14__9__sv2v_reg ,\xz.mem_with_zero_14__8__sv2v_reg ,
  \xz.mem_with_zero_14__7__sv2v_reg ,\xz.mem_with_zero_14__6__sv2v_reg ,
  \xz.mem_with_zero_14__5__sv2v_reg ,\xz.mem_with_zero_14__4__sv2v_reg ,
  \xz.mem_with_zero_14__3__sv2v_reg ,\xz.mem_with_zero_14__2__sv2v_reg ,
  \xz.mem_with_zero_14__1__sv2v_reg ,\xz.mem_with_zero_14__0__sv2v_reg ,\xz.mem_with_zero_13__31__sv2v_reg ,
  \xz.mem_with_zero_13__30__sv2v_reg ,\xz.mem_with_zero_13__29__sv2v_reg ,
  \xz.mem_with_zero_13__28__sv2v_reg ,\xz.mem_with_zero_13__27__sv2v_reg ,
  \xz.mem_with_zero_13__26__sv2v_reg ,\xz.mem_with_zero_13__25__sv2v_reg ,
  \xz.mem_with_zero_13__24__sv2v_reg ,\xz.mem_with_zero_13__23__sv2v_reg ,\xz.mem_with_zero_13__22__sv2v_reg ,
  \xz.mem_with_zero_13__21__sv2v_reg ,\xz.mem_with_zero_13__20__sv2v_reg ,
  \xz.mem_with_zero_13__19__sv2v_reg ,\xz.mem_with_zero_13__18__sv2v_reg ,
  \xz.mem_with_zero_13__17__sv2v_reg ,\xz.mem_with_zero_13__16__sv2v_reg ,
  \xz.mem_with_zero_13__15__sv2v_reg ,\xz.mem_with_zero_13__14__sv2v_reg ,\xz.mem_with_zero_13__13__sv2v_reg ,
  \xz.mem_with_zero_13__12__sv2v_reg ,\xz.mem_with_zero_13__11__sv2v_reg ,
  \xz.mem_with_zero_13__10__sv2v_reg ,\xz.mem_with_zero_13__9__sv2v_reg ,
  \xz.mem_with_zero_13__8__sv2v_reg ,\xz.mem_with_zero_13__7__sv2v_reg ,
  \xz.mem_with_zero_13__6__sv2v_reg ,\xz.mem_with_zero_13__5__sv2v_reg ,\xz.mem_with_zero_13__4__sv2v_reg ,
  \xz.mem_with_zero_13__3__sv2v_reg ,\xz.mem_with_zero_13__2__sv2v_reg ,
  \xz.mem_with_zero_13__1__sv2v_reg ,\xz.mem_with_zero_13__0__sv2v_reg ,
  \xz.mem_with_zero_12__31__sv2v_reg ,\xz.mem_with_zero_12__30__sv2v_reg ,
  \xz.mem_with_zero_12__29__sv2v_reg ,\xz.mem_with_zero_12__28__sv2v_reg ,\xz.mem_with_zero_12__27__sv2v_reg ,
  \xz.mem_with_zero_12__26__sv2v_reg ,\xz.mem_with_zero_12__25__sv2v_reg ,
  \xz.mem_with_zero_12__24__sv2v_reg ,\xz.mem_with_zero_12__23__sv2v_reg ,
  \xz.mem_with_zero_12__22__sv2v_reg ,\xz.mem_with_zero_12__21__sv2v_reg ,
  \xz.mem_with_zero_12__20__sv2v_reg ,\xz.mem_with_zero_12__19__sv2v_reg ,
  \xz.mem_with_zero_12__18__sv2v_reg ,\xz.mem_with_zero_12__17__sv2v_reg ,\xz.mem_with_zero_12__16__sv2v_reg ,
  \xz.mem_with_zero_12__15__sv2v_reg ,\xz.mem_with_zero_12__14__sv2v_reg ,
  \xz.mem_with_zero_12__13__sv2v_reg ,\xz.mem_with_zero_12__12__sv2v_reg ,
  \xz.mem_with_zero_12__11__sv2v_reg ,\xz.mem_with_zero_12__10__sv2v_reg ,
  \xz.mem_with_zero_12__9__sv2v_reg ,\xz.mem_with_zero_12__8__sv2v_reg ,\xz.mem_with_zero_12__7__sv2v_reg ,
  \xz.mem_with_zero_12__6__sv2v_reg ,\xz.mem_with_zero_12__5__sv2v_reg ,
  \xz.mem_with_zero_12__4__sv2v_reg ,\xz.mem_with_zero_12__3__sv2v_reg ,
  \xz.mem_with_zero_12__2__sv2v_reg ,\xz.mem_with_zero_12__1__sv2v_reg ,\xz.mem_with_zero_12__0__sv2v_reg ,
  \xz.mem_with_zero_11__31__sv2v_reg ,\xz.mem_with_zero_11__30__sv2v_reg ,
  \xz.mem_with_zero_11__29__sv2v_reg ,\xz.mem_with_zero_11__28__sv2v_reg ,
  \xz.mem_with_zero_11__27__sv2v_reg ,\xz.mem_with_zero_11__26__sv2v_reg ,
  \xz.mem_with_zero_11__25__sv2v_reg ,\xz.mem_with_zero_11__24__sv2v_reg ,
  \xz.mem_with_zero_11__23__sv2v_reg ,\xz.mem_with_zero_11__22__sv2v_reg ,\xz.mem_with_zero_11__21__sv2v_reg ,
  \xz.mem_with_zero_11__20__sv2v_reg ,\xz.mem_with_zero_11__19__sv2v_reg ,
  \xz.mem_with_zero_11__18__sv2v_reg ,\xz.mem_with_zero_11__17__sv2v_reg ,
  \xz.mem_with_zero_11__16__sv2v_reg ,\xz.mem_with_zero_11__15__sv2v_reg ,
  \xz.mem_with_zero_11__14__sv2v_reg ,\xz.mem_with_zero_11__13__sv2v_reg ,\xz.mem_with_zero_11__12__sv2v_reg ,
  \xz.mem_with_zero_11__11__sv2v_reg ,\xz.mem_with_zero_11__10__sv2v_reg ,
  \xz.mem_with_zero_11__9__sv2v_reg ,\xz.mem_with_zero_11__8__sv2v_reg ,
  \xz.mem_with_zero_11__7__sv2v_reg ,\xz.mem_with_zero_11__6__sv2v_reg ,
  \xz.mem_with_zero_11__5__sv2v_reg ,\xz.mem_with_zero_11__4__sv2v_reg ,\xz.mem_with_zero_11__3__sv2v_reg ,
  \xz.mem_with_zero_11__2__sv2v_reg ,\xz.mem_with_zero_11__1__sv2v_reg ,
  \xz.mem_with_zero_11__0__sv2v_reg ,\xz.mem_with_zero_10__31__sv2v_reg ,
  \xz.mem_with_zero_10__30__sv2v_reg ,\xz.mem_with_zero_10__29__sv2v_reg ,
  \xz.mem_with_zero_10__28__sv2v_reg ,\xz.mem_with_zero_10__27__sv2v_reg ,\xz.mem_with_zero_10__26__sv2v_reg ,
  \xz.mem_with_zero_10__25__sv2v_reg ,\xz.mem_with_zero_10__24__sv2v_reg ,
  \xz.mem_with_zero_10__23__sv2v_reg ,\xz.mem_with_zero_10__22__sv2v_reg ,
  \xz.mem_with_zero_10__21__sv2v_reg ,\xz.mem_with_zero_10__20__sv2v_reg ,
  \xz.mem_with_zero_10__19__sv2v_reg ,\xz.mem_with_zero_10__18__sv2v_reg ,
  \xz.mem_with_zero_10__17__sv2v_reg ,\xz.mem_with_zero_10__16__sv2v_reg ,\xz.mem_with_zero_10__15__sv2v_reg ,
  \xz.mem_with_zero_10__14__sv2v_reg ,\xz.mem_with_zero_10__13__sv2v_reg ,
  \xz.mem_with_zero_10__12__sv2v_reg ,\xz.mem_with_zero_10__11__sv2v_reg ,
  \xz.mem_with_zero_10__10__sv2v_reg ,\xz.mem_with_zero_10__9__sv2v_reg ,
  \xz.mem_with_zero_10__8__sv2v_reg ,\xz.mem_with_zero_10__7__sv2v_reg ,\xz.mem_with_zero_10__6__sv2v_reg ,
  \xz.mem_with_zero_10__5__sv2v_reg ,\xz.mem_with_zero_10__4__sv2v_reg ,
  \xz.mem_with_zero_10__3__sv2v_reg ,\xz.mem_with_zero_10__2__sv2v_reg ,
  \xz.mem_with_zero_10__1__sv2v_reg ,\xz.mem_with_zero_10__0__sv2v_reg ,\xz.mem_with_zero_9__31__sv2v_reg ,
  \xz.mem_with_zero_9__30__sv2v_reg ,\xz.mem_with_zero_9__29__sv2v_reg ,
  \xz.mem_with_zero_9__28__sv2v_reg ,\xz.mem_with_zero_9__27__sv2v_reg ,
  \xz.mem_with_zero_9__26__sv2v_reg ,\xz.mem_with_zero_9__25__sv2v_reg ,
  \xz.mem_with_zero_9__24__sv2v_reg ,\xz.mem_with_zero_9__23__sv2v_reg ,\xz.mem_with_zero_9__22__sv2v_reg ,
  \xz.mem_with_zero_9__21__sv2v_reg ,\xz.mem_with_zero_9__20__sv2v_reg ,
  \xz.mem_with_zero_9__19__sv2v_reg ,\xz.mem_with_zero_9__18__sv2v_reg ,
  \xz.mem_with_zero_9__17__sv2v_reg ,\xz.mem_with_zero_9__16__sv2v_reg ,\xz.mem_with_zero_9__15__sv2v_reg ,
  \xz.mem_with_zero_9__14__sv2v_reg ,\xz.mem_with_zero_9__13__sv2v_reg ,
  \xz.mem_with_zero_9__12__sv2v_reg ,\xz.mem_with_zero_9__11__sv2v_reg ,
  \xz.mem_with_zero_9__10__sv2v_reg ,\xz.mem_with_zero_9__9__sv2v_reg ,
  \xz.mem_with_zero_9__8__sv2v_reg ,\xz.mem_with_zero_9__7__sv2v_reg ,\xz.mem_with_zero_9__6__sv2v_reg ,
  \xz.mem_with_zero_9__5__sv2v_reg ,\xz.mem_with_zero_9__4__sv2v_reg ,
  \xz.mem_with_zero_9__3__sv2v_reg ,\xz.mem_with_zero_9__2__sv2v_reg ,\xz.mem_with_zero_9__1__sv2v_reg ,
  \xz.mem_with_zero_9__0__sv2v_reg ,\xz.mem_with_zero_8__31__sv2v_reg ,
  \xz.mem_with_zero_8__30__sv2v_reg ,\xz.mem_with_zero_8__29__sv2v_reg ,
  \xz.mem_with_zero_8__28__sv2v_reg ,\xz.mem_with_zero_8__27__sv2v_reg ,
  \xz.mem_with_zero_8__26__sv2v_reg ,\xz.mem_with_zero_8__25__sv2v_reg ,\xz.mem_with_zero_8__24__sv2v_reg ,
  \xz.mem_with_zero_8__23__sv2v_reg ,\xz.mem_with_zero_8__22__sv2v_reg ,
  \xz.mem_with_zero_8__21__sv2v_reg ,\xz.mem_with_zero_8__20__sv2v_reg ,
  \xz.mem_with_zero_8__19__sv2v_reg ,\xz.mem_with_zero_8__18__sv2v_reg ,\xz.mem_with_zero_8__17__sv2v_reg ,
  \xz.mem_with_zero_8__16__sv2v_reg ,\xz.mem_with_zero_8__15__sv2v_reg ,
  \xz.mem_with_zero_8__14__sv2v_reg ,\xz.mem_with_zero_8__13__sv2v_reg ,
  \xz.mem_with_zero_8__12__sv2v_reg ,\xz.mem_with_zero_8__11__sv2v_reg ,
  \xz.mem_with_zero_8__10__sv2v_reg ,\xz.mem_with_zero_8__9__sv2v_reg ,\xz.mem_with_zero_8__8__sv2v_reg ,
  \xz.mem_with_zero_8__7__sv2v_reg ,\xz.mem_with_zero_8__6__sv2v_reg ,
  \xz.mem_with_zero_8__5__sv2v_reg ,\xz.mem_with_zero_8__4__sv2v_reg ,
  \xz.mem_with_zero_8__3__sv2v_reg ,\xz.mem_with_zero_8__2__sv2v_reg ,\xz.mem_with_zero_8__1__sv2v_reg ,
  \xz.mem_with_zero_8__0__sv2v_reg ,\xz.mem_with_zero_7__31__sv2v_reg ,
  \xz.mem_with_zero_7__30__sv2v_reg ,\xz.mem_with_zero_7__29__sv2v_reg ,
  \xz.mem_with_zero_7__28__sv2v_reg ,\xz.mem_with_zero_7__27__sv2v_reg ,\xz.mem_with_zero_7__26__sv2v_reg ,
  \xz.mem_with_zero_7__25__sv2v_reg ,\xz.mem_with_zero_7__24__sv2v_reg ,
  \xz.mem_with_zero_7__23__sv2v_reg ,\xz.mem_with_zero_7__22__sv2v_reg ,
  \xz.mem_with_zero_7__21__sv2v_reg ,\xz.mem_with_zero_7__20__sv2v_reg ,\xz.mem_with_zero_7__19__sv2v_reg ,
  \xz.mem_with_zero_7__18__sv2v_reg ,\xz.mem_with_zero_7__17__sv2v_reg ,
  \xz.mem_with_zero_7__16__sv2v_reg ,\xz.mem_with_zero_7__15__sv2v_reg ,
  \xz.mem_with_zero_7__14__sv2v_reg ,\xz.mem_with_zero_7__13__sv2v_reg ,
  \xz.mem_with_zero_7__12__sv2v_reg ,\xz.mem_with_zero_7__11__sv2v_reg ,\xz.mem_with_zero_7__10__sv2v_reg ,
  \xz.mem_with_zero_7__9__sv2v_reg ,\xz.mem_with_zero_7__8__sv2v_reg ,
  \xz.mem_with_zero_7__7__sv2v_reg ,\xz.mem_with_zero_7__6__sv2v_reg ,
  \xz.mem_with_zero_7__5__sv2v_reg ,\xz.mem_with_zero_7__4__sv2v_reg ,\xz.mem_with_zero_7__3__sv2v_reg ,
  \xz.mem_with_zero_7__2__sv2v_reg ,\xz.mem_with_zero_7__1__sv2v_reg ,
  \xz.mem_with_zero_7__0__sv2v_reg ,\xz.mem_with_zero_6__31__sv2v_reg ,
  \xz.mem_with_zero_6__30__sv2v_reg ,\xz.mem_with_zero_6__29__sv2v_reg ,\xz.mem_with_zero_6__28__sv2v_reg ,
  \xz.mem_with_zero_6__27__sv2v_reg ,\xz.mem_with_zero_6__26__sv2v_reg ,
  \xz.mem_with_zero_6__25__sv2v_reg ,\xz.mem_with_zero_6__24__sv2v_reg ,
  \xz.mem_with_zero_6__23__sv2v_reg ,\xz.mem_with_zero_6__22__sv2v_reg ,\xz.mem_with_zero_6__21__sv2v_reg ,
  \xz.mem_with_zero_6__20__sv2v_reg ,\xz.mem_with_zero_6__19__sv2v_reg ,
  \xz.mem_with_zero_6__18__sv2v_reg ,\xz.mem_with_zero_6__17__sv2v_reg ,
  \xz.mem_with_zero_6__16__sv2v_reg ,\xz.mem_with_zero_6__15__sv2v_reg ,
  \xz.mem_with_zero_6__14__sv2v_reg ,\xz.mem_with_zero_6__13__sv2v_reg ,\xz.mem_with_zero_6__12__sv2v_reg ,
  \xz.mem_with_zero_6__11__sv2v_reg ,\xz.mem_with_zero_6__10__sv2v_reg ,
  \xz.mem_with_zero_6__9__sv2v_reg ,\xz.mem_with_zero_6__8__sv2v_reg ,
  \xz.mem_with_zero_6__7__sv2v_reg ,\xz.mem_with_zero_6__6__sv2v_reg ,\xz.mem_with_zero_6__5__sv2v_reg ,
  \xz.mem_with_zero_6__4__sv2v_reg ,\xz.mem_with_zero_6__3__sv2v_reg ,
  \xz.mem_with_zero_6__2__sv2v_reg ,\xz.mem_with_zero_6__1__sv2v_reg ,
  \xz.mem_with_zero_6__0__sv2v_reg ,\xz.mem_with_zero_5__31__sv2v_reg ,\xz.mem_with_zero_5__30__sv2v_reg ,
  \xz.mem_with_zero_5__29__sv2v_reg ,\xz.mem_with_zero_5__28__sv2v_reg ,
  \xz.mem_with_zero_5__27__sv2v_reg ,\xz.mem_with_zero_5__26__sv2v_reg ,
  \xz.mem_with_zero_5__25__sv2v_reg ,\xz.mem_with_zero_5__24__sv2v_reg ,\xz.mem_with_zero_5__23__sv2v_reg ,
  \xz.mem_with_zero_5__22__sv2v_reg ,\xz.mem_with_zero_5__21__sv2v_reg ,
  \xz.mem_with_zero_5__20__sv2v_reg ,\xz.mem_with_zero_5__19__sv2v_reg ,
  \xz.mem_with_zero_5__18__sv2v_reg ,\xz.mem_with_zero_5__17__sv2v_reg ,
  \xz.mem_with_zero_5__16__sv2v_reg ,\xz.mem_with_zero_5__15__sv2v_reg ,\xz.mem_with_zero_5__14__sv2v_reg ,
  \xz.mem_with_zero_5__13__sv2v_reg ,\xz.mem_with_zero_5__12__sv2v_reg ,
  \xz.mem_with_zero_5__11__sv2v_reg ,\xz.mem_with_zero_5__10__sv2v_reg ,
  \xz.mem_with_zero_5__9__sv2v_reg ,\xz.mem_with_zero_5__8__sv2v_reg ,\xz.mem_with_zero_5__7__sv2v_reg ,
  \xz.mem_with_zero_5__6__sv2v_reg ,\xz.mem_with_zero_5__5__sv2v_reg ,
  \xz.mem_with_zero_5__4__sv2v_reg ,\xz.mem_with_zero_5__3__sv2v_reg ,
  \xz.mem_with_zero_5__2__sv2v_reg ,\xz.mem_with_zero_5__1__sv2v_reg ,\xz.mem_with_zero_5__0__sv2v_reg ,
  \xz.mem_with_zero_4__31__sv2v_reg ,\xz.mem_with_zero_4__30__sv2v_reg ,
  \xz.mem_with_zero_4__29__sv2v_reg ,\xz.mem_with_zero_4__28__sv2v_reg ,
  \xz.mem_with_zero_4__27__sv2v_reg ,\xz.mem_with_zero_4__26__sv2v_reg ,\xz.mem_with_zero_4__25__sv2v_reg ,
  \xz.mem_with_zero_4__24__sv2v_reg ,\xz.mem_with_zero_4__23__sv2v_reg ,
  \xz.mem_with_zero_4__22__sv2v_reg ,\xz.mem_with_zero_4__21__sv2v_reg ,
  \xz.mem_with_zero_4__20__sv2v_reg ,\xz.mem_with_zero_4__19__sv2v_reg ,
  \xz.mem_with_zero_4__18__sv2v_reg ,\xz.mem_with_zero_4__17__sv2v_reg ,\xz.mem_with_zero_4__16__sv2v_reg ,
  \xz.mem_with_zero_4__15__sv2v_reg ,\xz.mem_with_zero_4__14__sv2v_reg ,
  \xz.mem_with_zero_4__13__sv2v_reg ,\xz.mem_with_zero_4__12__sv2v_reg ,
  \xz.mem_with_zero_4__11__sv2v_reg ,\xz.mem_with_zero_4__10__sv2v_reg ,\xz.mem_with_zero_4__9__sv2v_reg ,
  \xz.mem_with_zero_4__8__sv2v_reg ,\xz.mem_with_zero_4__7__sv2v_reg ,
  \xz.mem_with_zero_4__6__sv2v_reg ,\xz.mem_with_zero_4__5__sv2v_reg ,
  \xz.mem_with_zero_4__4__sv2v_reg ,\xz.mem_with_zero_4__3__sv2v_reg ,\xz.mem_with_zero_4__2__sv2v_reg ,
  \xz.mem_with_zero_4__1__sv2v_reg ,\xz.mem_with_zero_4__0__sv2v_reg ,
  \xz.mem_with_zero_3__31__sv2v_reg ,\xz.mem_with_zero_3__30__sv2v_reg ,
  \xz.mem_with_zero_3__29__sv2v_reg ,\xz.mem_with_zero_3__28__sv2v_reg ,\xz.mem_with_zero_3__27__sv2v_reg ,
  \xz.mem_with_zero_3__26__sv2v_reg ,\xz.mem_with_zero_3__25__sv2v_reg ,
  \xz.mem_with_zero_3__24__sv2v_reg ,\xz.mem_with_zero_3__23__sv2v_reg ,
  \xz.mem_with_zero_3__22__sv2v_reg ,\xz.mem_with_zero_3__21__sv2v_reg ,
  \xz.mem_with_zero_3__20__sv2v_reg ,\xz.mem_with_zero_3__19__sv2v_reg ,\xz.mem_with_zero_3__18__sv2v_reg ,
  \xz.mem_with_zero_3__17__sv2v_reg ,\xz.mem_with_zero_3__16__sv2v_reg ,
  \xz.mem_with_zero_3__15__sv2v_reg ,\xz.mem_with_zero_3__14__sv2v_reg ,
  \xz.mem_with_zero_3__13__sv2v_reg ,\xz.mem_with_zero_3__12__sv2v_reg ,\xz.mem_with_zero_3__11__sv2v_reg ,
  \xz.mem_with_zero_3__10__sv2v_reg ,\xz.mem_with_zero_3__9__sv2v_reg ,
  \xz.mem_with_zero_3__8__sv2v_reg ,\xz.mem_with_zero_3__7__sv2v_reg ,
  \xz.mem_with_zero_3__6__sv2v_reg ,\xz.mem_with_zero_3__5__sv2v_reg ,\xz.mem_with_zero_3__4__sv2v_reg ,
  \xz.mem_with_zero_3__3__sv2v_reg ,\xz.mem_with_zero_3__2__sv2v_reg ,
  \xz.mem_with_zero_3__1__sv2v_reg ,\xz.mem_with_zero_3__0__sv2v_reg ,
  \xz.mem_with_zero_2__31__sv2v_reg ,\xz.mem_with_zero_2__30__sv2v_reg ,\xz.mem_with_zero_2__29__sv2v_reg ,
  \xz.mem_with_zero_2__28__sv2v_reg ,\xz.mem_with_zero_2__27__sv2v_reg ,
  \xz.mem_with_zero_2__26__sv2v_reg ,\xz.mem_with_zero_2__25__sv2v_reg ,
  \xz.mem_with_zero_2__24__sv2v_reg ,\xz.mem_with_zero_2__23__sv2v_reg ,
  \xz.mem_with_zero_2__22__sv2v_reg ,\xz.mem_with_zero_2__21__sv2v_reg ,\xz.mem_with_zero_2__20__sv2v_reg ,
  \xz.mem_with_zero_2__19__sv2v_reg ,\xz.mem_with_zero_2__18__sv2v_reg ,
  \xz.mem_with_zero_2__17__sv2v_reg ,\xz.mem_with_zero_2__16__sv2v_reg ,
  \xz.mem_with_zero_2__15__sv2v_reg ,\xz.mem_with_zero_2__14__sv2v_reg ,\xz.mem_with_zero_2__13__sv2v_reg ,
  \xz.mem_with_zero_2__12__sv2v_reg ,\xz.mem_with_zero_2__11__sv2v_reg ,
  \xz.mem_with_zero_2__10__sv2v_reg ,\xz.mem_with_zero_2__9__sv2v_reg ,
  \xz.mem_with_zero_2__8__sv2v_reg ,\xz.mem_with_zero_2__7__sv2v_reg ,\xz.mem_with_zero_2__6__sv2v_reg ,
  \xz.mem_with_zero_2__5__sv2v_reg ,\xz.mem_with_zero_2__4__sv2v_reg ,
  \xz.mem_with_zero_2__3__sv2v_reg ,\xz.mem_with_zero_2__2__sv2v_reg ,
  \xz.mem_with_zero_2__1__sv2v_reg ,\xz.mem_with_zero_2__0__sv2v_reg ,\xz.mem_with_zero_1__31__sv2v_reg ,
  \xz.mem_with_zero_1__30__sv2v_reg ,\xz.mem_with_zero_1__29__sv2v_reg ,
  \xz.mem_with_zero_1__28__sv2v_reg ,\xz.mem_with_zero_1__27__sv2v_reg ,
  \xz.mem_with_zero_1__26__sv2v_reg ,\xz.mem_with_zero_1__25__sv2v_reg ,
  \xz.mem_with_zero_1__24__sv2v_reg ,\xz.mem_with_zero_1__23__sv2v_reg ,\xz.mem_with_zero_1__22__sv2v_reg ,
  \xz.mem_with_zero_1__21__sv2v_reg ,\xz.mem_with_zero_1__20__sv2v_reg ,
  \xz.mem_with_zero_1__19__sv2v_reg ,\xz.mem_with_zero_1__18__sv2v_reg ,
  \xz.mem_with_zero_1__17__sv2v_reg ,\xz.mem_with_zero_1__16__sv2v_reg ,\xz.mem_with_zero_1__15__sv2v_reg ,
  \xz.mem_with_zero_1__14__sv2v_reg ,\xz.mem_with_zero_1__13__sv2v_reg ,
  \xz.mem_with_zero_1__12__sv2v_reg ,\xz.mem_with_zero_1__11__sv2v_reg ,
  \xz.mem_with_zero_1__10__sv2v_reg ,\xz.mem_with_zero_1__9__sv2v_reg ,
  \xz.mem_with_zero_1__8__sv2v_reg ,\xz.mem_with_zero_1__7__sv2v_reg ,\xz.mem_with_zero_1__6__sv2v_reg ,
  \xz.mem_with_zero_1__5__sv2v_reg ,\xz.mem_with_zero_1__4__sv2v_reg ,
  \xz.mem_with_zero_1__3__sv2v_reg ,\xz.mem_with_zero_1__2__sv2v_reg ,\xz.mem_with_zero_1__1__sv2v_reg ,
  \xz.mem_with_zero_1__0__sv2v_reg ;
  assign r_addr_r[9] = r_addr_r_9_sv2v_reg;
  assign r_addr_r[8] = r_addr_r_8_sv2v_reg;
  assign r_addr_r[7] = r_addr_r_7_sv2v_reg;
  assign r_addr_r[6] = r_addr_r_6_sv2v_reg;
  assign r_addr_r[5] = r_addr_r_5_sv2v_reg;
  assign r_addr_r[4] = r_addr_r_4_sv2v_reg;
  assign r_addr_r[3] = r_addr_r_3_sv2v_reg;
  assign r_addr_r[2] = r_addr_r_2_sv2v_reg;
  assign r_addr_r[1] = r_addr_r_1_sv2v_reg;
  assign r_addr_r[0] = r_addr_r_0_sv2v_reg;
  assign \xz.mem_with_zero_31__31_  = \xz.mem_with_zero_31__31__sv2v_reg ;
  assign \xz.mem_with_zero_31__30_  = \xz.mem_with_zero_31__30__sv2v_reg ;
  assign \xz.mem_with_zero_31__29_  = \xz.mem_with_zero_31__29__sv2v_reg ;
  assign \xz.mem_with_zero_31__28_  = \xz.mem_with_zero_31__28__sv2v_reg ;
  assign \xz.mem_with_zero_31__27_  = \xz.mem_with_zero_31__27__sv2v_reg ;
  assign \xz.mem_with_zero_31__26_  = \xz.mem_with_zero_31__26__sv2v_reg ;
  assign \xz.mem_with_zero_31__25_  = \xz.mem_with_zero_31__25__sv2v_reg ;
  assign \xz.mem_with_zero_31__24_  = \xz.mem_with_zero_31__24__sv2v_reg ;
  assign \xz.mem_with_zero_31__23_  = \xz.mem_with_zero_31__23__sv2v_reg ;
  assign \xz.mem_with_zero_31__22_  = \xz.mem_with_zero_31__22__sv2v_reg ;
  assign \xz.mem_with_zero_31__21_  = \xz.mem_with_zero_31__21__sv2v_reg ;
  assign \xz.mem_with_zero_31__20_  = \xz.mem_with_zero_31__20__sv2v_reg ;
  assign \xz.mem_with_zero_31__19_  = \xz.mem_with_zero_31__19__sv2v_reg ;
  assign \xz.mem_with_zero_31__18_  = \xz.mem_with_zero_31__18__sv2v_reg ;
  assign \xz.mem_with_zero_31__17_  = \xz.mem_with_zero_31__17__sv2v_reg ;
  assign \xz.mem_with_zero_31__16_  = \xz.mem_with_zero_31__16__sv2v_reg ;
  assign \xz.mem_with_zero_31__15_  = \xz.mem_with_zero_31__15__sv2v_reg ;
  assign \xz.mem_with_zero_31__14_  = \xz.mem_with_zero_31__14__sv2v_reg ;
  assign \xz.mem_with_zero_31__13_  = \xz.mem_with_zero_31__13__sv2v_reg ;
  assign \xz.mem_with_zero_31__12_  = \xz.mem_with_zero_31__12__sv2v_reg ;
  assign \xz.mem_with_zero_31__11_  = \xz.mem_with_zero_31__11__sv2v_reg ;
  assign \xz.mem_with_zero_31__10_  = \xz.mem_with_zero_31__10__sv2v_reg ;
  assign \xz.mem_with_zero_31__9_  = \xz.mem_with_zero_31__9__sv2v_reg ;
  assign \xz.mem_with_zero_31__8_  = \xz.mem_with_zero_31__8__sv2v_reg ;
  assign \xz.mem_with_zero_31__7_  = \xz.mem_with_zero_31__7__sv2v_reg ;
  assign \xz.mem_with_zero_31__6_  = \xz.mem_with_zero_31__6__sv2v_reg ;
  assign \xz.mem_with_zero_31__5_  = \xz.mem_with_zero_31__5__sv2v_reg ;
  assign \xz.mem_with_zero_31__4_  = \xz.mem_with_zero_31__4__sv2v_reg ;
  assign \xz.mem_with_zero_31__3_  = \xz.mem_with_zero_31__3__sv2v_reg ;
  assign \xz.mem_with_zero_31__2_  = \xz.mem_with_zero_31__2__sv2v_reg ;
  assign \xz.mem_with_zero_31__1_  = \xz.mem_with_zero_31__1__sv2v_reg ;
  assign \xz.mem_with_zero_31__0_  = \xz.mem_with_zero_31__0__sv2v_reg ;
  assign \xz.mem_with_zero_30__31_  = \xz.mem_with_zero_30__31__sv2v_reg ;
  assign \xz.mem_with_zero_30__30_  = \xz.mem_with_zero_30__30__sv2v_reg ;
  assign \xz.mem_with_zero_30__29_  = \xz.mem_with_zero_30__29__sv2v_reg ;
  assign \xz.mem_with_zero_30__28_  = \xz.mem_with_zero_30__28__sv2v_reg ;
  assign \xz.mem_with_zero_30__27_  = \xz.mem_with_zero_30__27__sv2v_reg ;
  assign \xz.mem_with_zero_30__26_  = \xz.mem_with_zero_30__26__sv2v_reg ;
  assign \xz.mem_with_zero_30__25_  = \xz.mem_with_zero_30__25__sv2v_reg ;
  assign \xz.mem_with_zero_30__24_  = \xz.mem_with_zero_30__24__sv2v_reg ;
  assign \xz.mem_with_zero_30__23_  = \xz.mem_with_zero_30__23__sv2v_reg ;
  assign \xz.mem_with_zero_30__22_  = \xz.mem_with_zero_30__22__sv2v_reg ;
  assign \xz.mem_with_zero_30__21_  = \xz.mem_with_zero_30__21__sv2v_reg ;
  assign \xz.mem_with_zero_30__20_  = \xz.mem_with_zero_30__20__sv2v_reg ;
  assign \xz.mem_with_zero_30__19_  = \xz.mem_with_zero_30__19__sv2v_reg ;
  assign \xz.mem_with_zero_30__18_  = \xz.mem_with_zero_30__18__sv2v_reg ;
  assign \xz.mem_with_zero_30__17_  = \xz.mem_with_zero_30__17__sv2v_reg ;
  assign \xz.mem_with_zero_30__16_  = \xz.mem_with_zero_30__16__sv2v_reg ;
  assign \xz.mem_with_zero_30__15_  = \xz.mem_with_zero_30__15__sv2v_reg ;
  assign \xz.mem_with_zero_30__14_  = \xz.mem_with_zero_30__14__sv2v_reg ;
  assign \xz.mem_with_zero_30__13_  = \xz.mem_with_zero_30__13__sv2v_reg ;
  assign \xz.mem_with_zero_30__12_  = \xz.mem_with_zero_30__12__sv2v_reg ;
  assign \xz.mem_with_zero_30__11_  = \xz.mem_with_zero_30__11__sv2v_reg ;
  assign \xz.mem_with_zero_30__10_  = \xz.mem_with_zero_30__10__sv2v_reg ;
  assign \xz.mem_with_zero_30__9_  = \xz.mem_with_zero_30__9__sv2v_reg ;
  assign \xz.mem_with_zero_30__8_  = \xz.mem_with_zero_30__8__sv2v_reg ;
  assign \xz.mem_with_zero_30__7_  = \xz.mem_with_zero_30__7__sv2v_reg ;
  assign \xz.mem_with_zero_30__6_  = \xz.mem_with_zero_30__6__sv2v_reg ;
  assign \xz.mem_with_zero_30__5_  = \xz.mem_with_zero_30__5__sv2v_reg ;
  assign \xz.mem_with_zero_30__4_  = \xz.mem_with_zero_30__4__sv2v_reg ;
  assign \xz.mem_with_zero_30__3_  = \xz.mem_with_zero_30__3__sv2v_reg ;
  assign \xz.mem_with_zero_30__2_  = \xz.mem_with_zero_30__2__sv2v_reg ;
  assign \xz.mem_with_zero_30__1_  = \xz.mem_with_zero_30__1__sv2v_reg ;
  assign \xz.mem_with_zero_30__0_  = \xz.mem_with_zero_30__0__sv2v_reg ;
  assign \xz.mem_with_zero_29__31_  = \xz.mem_with_zero_29__31__sv2v_reg ;
  assign \xz.mem_with_zero_29__30_  = \xz.mem_with_zero_29__30__sv2v_reg ;
  assign \xz.mem_with_zero_29__29_  = \xz.mem_with_zero_29__29__sv2v_reg ;
  assign \xz.mem_with_zero_29__28_  = \xz.mem_with_zero_29__28__sv2v_reg ;
  assign \xz.mem_with_zero_29__27_  = \xz.mem_with_zero_29__27__sv2v_reg ;
  assign \xz.mem_with_zero_29__26_  = \xz.mem_with_zero_29__26__sv2v_reg ;
  assign \xz.mem_with_zero_29__25_  = \xz.mem_with_zero_29__25__sv2v_reg ;
  assign \xz.mem_with_zero_29__24_  = \xz.mem_with_zero_29__24__sv2v_reg ;
  assign \xz.mem_with_zero_29__23_  = \xz.mem_with_zero_29__23__sv2v_reg ;
  assign \xz.mem_with_zero_29__22_  = \xz.mem_with_zero_29__22__sv2v_reg ;
  assign \xz.mem_with_zero_29__21_  = \xz.mem_with_zero_29__21__sv2v_reg ;
  assign \xz.mem_with_zero_29__20_  = \xz.mem_with_zero_29__20__sv2v_reg ;
  assign \xz.mem_with_zero_29__19_  = \xz.mem_with_zero_29__19__sv2v_reg ;
  assign \xz.mem_with_zero_29__18_  = \xz.mem_with_zero_29__18__sv2v_reg ;
  assign \xz.mem_with_zero_29__17_  = \xz.mem_with_zero_29__17__sv2v_reg ;
  assign \xz.mem_with_zero_29__16_  = \xz.mem_with_zero_29__16__sv2v_reg ;
  assign \xz.mem_with_zero_29__15_  = \xz.mem_with_zero_29__15__sv2v_reg ;
  assign \xz.mem_with_zero_29__14_  = \xz.mem_with_zero_29__14__sv2v_reg ;
  assign \xz.mem_with_zero_29__13_  = \xz.mem_with_zero_29__13__sv2v_reg ;
  assign \xz.mem_with_zero_29__12_  = \xz.mem_with_zero_29__12__sv2v_reg ;
  assign \xz.mem_with_zero_29__11_  = \xz.mem_with_zero_29__11__sv2v_reg ;
  assign \xz.mem_with_zero_29__10_  = \xz.mem_with_zero_29__10__sv2v_reg ;
  assign \xz.mem_with_zero_29__9_  = \xz.mem_with_zero_29__9__sv2v_reg ;
  assign \xz.mem_with_zero_29__8_  = \xz.mem_with_zero_29__8__sv2v_reg ;
  assign \xz.mem_with_zero_29__7_  = \xz.mem_with_zero_29__7__sv2v_reg ;
  assign \xz.mem_with_zero_29__6_  = \xz.mem_with_zero_29__6__sv2v_reg ;
  assign \xz.mem_with_zero_29__5_  = \xz.mem_with_zero_29__5__sv2v_reg ;
  assign \xz.mem_with_zero_29__4_  = \xz.mem_with_zero_29__4__sv2v_reg ;
  assign \xz.mem_with_zero_29__3_  = \xz.mem_with_zero_29__3__sv2v_reg ;
  assign \xz.mem_with_zero_29__2_  = \xz.mem_with_zero_29__2__sv2v_reg ;
  assign \xz.mem_with_zero_29__1_  = \xz.mem_with_zero_29__1__sv2v_reg ;
  assign \xz.mem_with_zero_29__0_  = \xz.mem_with_zero_29__0__sv2v_reg ;
  assign \xz.mem_with_zero_28__31_  = \xz.mem_with_zero_28__31__sv2v_reg ;
  assign \xz.mem_with_zero_28__30_  = \xz.mem_with_zero_28__30__sv2v_reg ;
  assign \xz.mem_with_zero_28__29_  = \xz.mem_with_zero_28__29__sv2v_reg ;
  assign \xz.mem_with_zero_28__28_  = \xz.mem_with_zero_28__28__sv2v_reg ;
  assign \xz.mem_with_zero_28__27_  = \xz.mem_with_zero_28__27__sv2v_reg ;
  assign \xz.mem_with_zero_28__26_  = \xz.mem_with_zero_28__26__sv2v_reg ;
  assign \xz.mem_with_zero_28__25_  = \xz.mem_with_zero_28__25__sv2v_reg ;
  assign \xz.mem_with_zero_28__24_  = \xz.mem_with_zero_28__24__sv2v_reg ;
  assign \xz.mem_with_zero_28__23_  = \xz.mem_with_zero_28__23__sv2v_reg ;
  assign \xz.mem_with_zero_28__22_  = \xz.mem_with_zero_28__22__sv2v_reg ;
  assign \xz.mem_with_zero_28__21_  = \xz.mem_with_zero_28__21__sv2v_reg ;
  assign \xz.mem_with_zero_28__20_  = \xz.mem_with_zero_28__20__sv2v_reg ;
  assign \xz.mem_with_zero_28__19_  = \xz.mem_with_zero_28__19__sv2v_reg ;
  assign \xz.mem_with_zero_28__18_  = \xz.mem_with_zero_28__18__sv2v_reg ;
  assign \xz.mem_with_zero_28__17_  = \xz.mem_with_zero_28__17__sv2v_reg ;
  assign \xz.mem_with_zero_28__16_  = \xz.mem_with_zero_28__16__sv2v_reg ;
  assign \xz.mem_with_zero_28__15_  = \xz.mem_with_zero_28__15__sv2v_reg ;
  assign \xz.mem_with_zero_28__14_  = \xz.mem_with_zero_28__14__sv2v_reg ;
  assign \xz.mem_with_zero_28__13_  = \xz.mem_with_zero_28__13__sv2v_reg ;
  assign \xz.mem_with_zero_28__12_  = \xz.mem_with_zero_28__12__sv2v_reg ;
  assign \xz.mem_with_zero_28__11_  = \xz.mem_with_zero_28__11__sv2v_reg ;
  assign \xz.mem_with_zero_28__10_  = \xz.mem_with_zero_28__10__sv2v_reg ;
  assign \xz.mem_with_zero_28__9_  = \xz.mem_with_zero_28__9__sv2v_reg ;
  assign \xz.mem_with_zero_28__8_  = \xz.mem_with_zero_28__8__sv2v_reg ;
  assign \xz.mem_with_zero_28__7_  = \xz.mem_with_zero_28__7__sv2v_reg ;
  assign \xz.mem_with_zero_28__6_  = \xz.mem_with_zero_28__6__sv2v_reg ;
  assign \xz.mem_with_zero_28__5_  = \xz.mem_with_zero_28__5__sv2v_reg ;
  assign \xz.mem_with_zero_28__4_  = \xz.mem_with_zero_28__4__sv2v_reg ;
  assign \xz.mem_with_zero_28__3_  = \xz.mem_with_zero_28__3__sv2v_reg ;
  assign \xz.mem_with_zero_28__2_  = \xz.mem_with_zero_28__2__sv2v_reg ;
  assign \xz.mem_with_zero_28__1_  = \xz.mem_with_zero_28__1__sv2v_reg ;
  assign \xz.mem_with_zero_28__0_  = \xz.mem_with_zero_28__0__sv2v_reg ;
  assign \xz.mem_with_zero_27__31_  = \xz.mem_with_zero_27__31__sv2v_reg ;
  assign \xz.mem_with_zero_27__30_  = \xz.mem_with_zero_27__30__sv2v_reg ;
  assign \xz.mem_with_zero_27__29_  = \xz.mem_with_zero_27__29__sv2v_reg ;
  assign \xz.mem_with_zero_27__28_  = \xz.mem_with_zero_27__28__sv2v_reg ;
  assign \xz.mem_with_zero_27__27_  = \xz.mem_with_zero_27__27__sv2v_reg ;
  assign \xz.mem_with_zero_27__26_  = \xz.mem_with_zero_27__26__sv2v_reg ;
  assign \xz.mem_with_zero_27__25_  = \xz.mem_with_zero_27__25__sv2v_reg ;
  assign \xz.mem_with_zero_27__24_  = \xz.mem_with_zero_27__24__sv2v_reg ;
  assign \xz.mem_with_zero_27__23_  = \xz.mem_with_zero_27__23__sv2v_reg ;
  assign \xz.mem_with_zero_27__22_  = \xz.mem_with_zero_27__22__sv2v_reg ;
  assign \xz.mem_with_zero_27__21_  = \xz.mem_with_zero_27__21__sv2v_reg ;
  assign \xz.mem_with_zero_27__20_  = \xz.mem_with_zero_27__20__sv2v_reg ;
  assign \xz.mem_with_zero_27__19_  = \xz.mem_with_zero_27__19__sv2v_reg ;
  assign \xz.mem_with_zero_27__18_  = \xz.mem_with_zero_27__18__sv2v_reg ;
  assign \xz.mem_with_zero_27__17_  = \xz.mem_with_zero_27__17__sv2v_reg ;
  assign \xz.mem_with_zero_27__16_  = \xz.mem_with_zero_27__16__sv2v_reg ;
  assign \xz.mem_with_zero_27__15_  = \xz.mem_with_zero_27__15__sv2v_reg ;
  assign \xz.mem_with_zero_27__14_  = \xz.mem_with_zero_27__14__sv2v_reg ;
  assign \xz.mem_with_zero_27__13_  = \xz.mem_with_zero_27__13__sv2v_reg ;
  assign \xz.mem_with_zero_27__12_  = \xz.mem_with_zero_27__12__sv2v_reg ;
  assign \xz.mem_with_zero_27__11_  = \xz.mem_with_zero_27__11__sv2v_reg ;
  assign \xz.mem_with_zero_27__10_  = \xz.mem_with_zero_27__10__sv2v_reg ;
  assign \xz.mem_with_zero_27__9_  = \xz.mem_with_zero_27__9__sv2v_reg ;
  assign \xz.mem_with_zero_27__8_  = \xz.mem_with_zero_27__8__sv2v_reg ;
  assign \xz.mem_with_zero_27__7_  = \xz.mem_with_zero_27__7__sv2v_reg ;
  assign \xz.mem_with_zero_27__6_  = \xz.mem_with_zero_27__6__sv2v_reg ;
  assign \xz.mem_with_zero_27__5_  = \xz.mem_with_zero_27__5__sv2v_reg ;
  assign \xz.mem_with_zero_27__4_  = \xz.mem_with_zero_27__4__sv2v_reg ;
  assign \xz.mem_with_zero_27__3_  = \xz.mem_with_zero_27__3__sv2v_reg ;
  assign \xz.mem_with_zero_27__2_  = \xz.mem_with_zero_27__2__sv2v_reg ;
  assign \xz.mem_with_zero_27__1_  = \xz.mem_with_zero_27__1__sv2v_reg ;
  assign \xz.mem_with_zero_27__0_  = \xz.mem_with_zero_27__0__sv2v_reg ;
  assign \xz.mem_with_zero_26__31_  = \xz.mem_with_zero_26__31__sv2v_reg ;
  assign \xz.mem_with_zero_26__30_  = \xz.mem_with_zero_26__30__sv2v_reg ;
  assign \xz.mem_with_zero_26__29_  = \xz.mem_with_zero_26__29__sv2v_reg ;
  assign \xz.mem_with_zero_26__28_  = \xz.mem_with_zero_26__28__sv2v_reg ;
  assign \xz.mem_with_zero_26__27_  = \xz.mem_with_zero_26__27__sv2v_reg ;
  assign \xz.mem_with_zero_26__26_  = \xz.mem_with_zero_26__26__sv2v_reg ;
  assign \xz.mem_with_zero_26__25_  = \xz.mem_with_zero_26__25__sv2v_reg ;
  assign \xz.mem_with_zero_26__24_  = \xz.mem_with_zero_26__24__sv2v_reg ;
  assign \xz.mem_with_zero_26__23_  = \xz.mem_with_zero_26__23__sv2v_reg ;
  assign \xz.mem_with_zero_26__22_  = \xz.mem_with_zero_26__22__sv2v_reg ;
  assign \xz.mem_with_zero_26__21_  = \xz.mem_with_zero_26__21__sv2v_reg ;
  assign \xz.mem_with_zero_26__20_  = \xz.mem_with_zero_26__20__sv2v_reg ;
  assign \xz.mem_with_zero_26__19_  = \xz.mem_with_zero_26__19__sv2v_reg ;
  assign \xz.mem_with_zero_26__18_  = \xz.mem_with_zero_26__18__sv2v_reg ;
  assign \xz.mem_with_zero_26__17_  = \xz.mem_with_zero_26__17__sv2v_reg ;
  assign \xz.mem_with_zero_26__16_  = \xz.mem_with_zero_26__16__sv2v_reg ;
  assign \xz.mem_with_zero_26__15_  = \xz.mem_with_zero_26__15__sv2v_reg ;
  assign \xz.mem_with_zero_26__14_  = \xz.mem_with_zero_26__14__sv2v_reg ;
  assign \xz.mem_with_zero_26__13_  = \xz.mem_with_zero_26__13__sv2v_reg ;
  assign \xz.mem_with_zero_26__12_  = \xz.mem_with_zero_26__12__sv2v_reg ;
  assign \xz.mem_with_zero_26__11_  = \xz.mem_with_zero_26__11__sv2v_reg ;
  assign \xz.mem_with_zero_26__10_  = \xz.mem_with_zero_26__10__sv2v_reg ;
  assign \xz.mem_with_zero_26__9_  = \xz.mem_with_zero_26__9__sv2v_reg ;
  assign \xz.mem_with_zero_26__8_  = \xz.mem_with_zero_26__8__sv2v_reg ;
  assign \xz.mem_with_zero_26__7_  = \xz.mem_with_zero_26__7__sv2v_reg ;
  assign \xz.mem_with_zero_26__6_  = \xz.mem_with_zero_26__6__sv2v_reg ;
  assign \xz.mem_with_zero_26__5_  = \xz.mem_with_zero_26__5__sv2v_reg ;
  assign \xz.mem_with_zero_26__4_  = \xz.mem_with_zero_26__4__sv2v_reg ;
  assign \xz.mem_with_zero_26__3_  = \xz.mem_with_zero_26__3__sv2v_reg ;
  assign \xz.mem_with_zero_26__2_  = \xz.mem_with_zero_26__2__sv2v_reg ;
  assign \xz.mem_with_zero_26__1_  = \xz.mem_with_zero_26__1__sv2v_reg ;
  assign \xz.mem_with_zero_26__0_  = \xz.mem_with_zero_26__0__sv2v_reg ;
  assign \xz.mem_with_zero_25__31_  = \xz.mem_with_zero_25__31__sv2v_reg ;
  assign \xz.mem_with_zero_25__30_  = \xz.mem_with_zero_25__30__sv2v_reg ;
  assign \xz.mem_with_zero_25__29_  = \xz.mem_with_zero_25__29__sv2v_reg ;
  assign \xz.mem_with_zero_25__28_  = \xz.mem_with_zero_25__28__sv2v_reg ;
  assign \xz.mem_with_zero_25__27_  = \xz.mem_with_zero_25__27__sv2v_reg ;
  assign \xz.mem_with_zero_25__26_  = \xz.mem_with_zero_25__26__sv2v_reg ;
  assign \xz.mem_with_zero_25__25_  = \xz.mem_with_zero_25__25__sv2v_reg ;
  assign \xz.mem_with_zero_25__24_  = \xz.mem_with_zero_25__24__sv2v_reg ;
  assign \xz.mem_with_zero_25__23_  = \xz.mem_with_zero_25__23__sv2v_reg ;
  assign \xz.mem_with_zero_25__22_  = \xz.mem_with_zero_25__22__sv2v_reg ;
  assign \xz.mem_with_zero_25__21_  = \xz.mem_with_zero_25__21__sv2v_reg ;
  assign \xz.mem_with_zero_25__20_  = \xz.mem_with_zero_25__20__sv2v_reg ;
  assign \xz.mem_with_zero_25__19_  = \xz.mem_with_zero_25__19__sv2v_reg ;
  assign \xz.mem_with_zero_25__18_  = \xz.mem_with_zero_25__18__sv2v_reg ;
  assign \xz.mem_with_zero_25__17_  = \xz.mem_with_zero_25__17__sv2v_reg ;
  assign \xz.mem_with_zero_25__16_  = \xz.mem_with_zero_25__16__sv2v_reg ;
  assign \xz.mem_with_zero_25__15_  = \xz.mem_with_zero_25__15__sv2v_reg ;
  assign \xz.mem_with_zero_25__14_  = \xz.mem_with_zero_25__14__sv2v_reg ;
  assign \xz.mem_with_zero_25__13_  = \xz.mem_with_zero_25__13__sv2v_reg ;
  assign \xz.mem_with_zero_25__12_  = \xz.mem_with_zero_25__12__sv2v_reg ;
  assign \xz.mem_with_zero_25__11_  = \xz.mem_with_zero_25__11__sv2v_reg ;
  assign \xz.mem_with_zero_25__10_  = \xz.mem_with_zero_25__10__sv2v_reg ;
  assign \xz.mem_with_zero_25__9_  = \xz.mem_with_zero_25__9__sv2v_reg ;
  assign \xz.mem_with_zero_25__8_  = \xz.mem_with_zero_25__8__sv2v_reg ;
  assign \xz.mem_with_zero_25__7_  = \xz.mem_with_zero_25__7__sv2v_reg ;
  assign \xz.mem_with_zero_25__6_  = \xz.mem_with_zero_25__6__sv2v_reg ;
  assign \xz.mem_with_zero_25__5_  = \xz.mem_with_zero_25__5__sv2v_reg ;
  assign \xz.mem_with_zero_25__4_  = \xz.mem_with_zero_25__4__sv2v_reg ;
  assign \xz.mem_with_zero_25__3_  = \xz.mem_with_zero_25__3__sv2v_reg ;
  assign \xz.mem_with_zero_25__2_  = \xz.mem_with_zero_25__2__sv2v_reg ;
  assign \xz.mem_with_zero_25__1_  = \xz.mem_with_zero_25__1__sv2v_reg ;
  assign \xz.mem_with_zero_25__0_  = \xz.mem_with_zero_25__0__sv2v_reg ;
  assign \xz.mem_with_zero_24__31_  = \xz.mem_with_zero_24__31__sv2v_reg ;
  assign \xz.mem_with_zero_24__30_  = \xz.mem_with_zero_24__30__sv2v_reg ;
  assign \xz.mem_with_zero_24__29_  = \xz.mem_with_zero_24__29__sv2v_reg ;
  assign \xz.mem_with_zero_24__28_  = \xz.mem_with_zero_24__28__sv2v_reg ;
  assign \xz.mem_with_zero_24__27_  = \xz.mem_with_zero_24__27__sv2v_reg ;
  assign \xz.mem_with_zero_24__26_  = \xz.mem_with_zero_24__26__sv2v_reg ;
  assign \xz.mem_with_zero_24__25_  = \xz.mem_with_zero_24__25__sv2v_reg ;
  assign \xz.mem_with_zero_24__24_  = \xz.mem_with_zero_24__24__sv2v_reg ;
  assign \xz.mem_with_zero_24__23_  = \xz.mem_with_zero_24__23__sv2v_reg ;
  assign \xz.mem_with_zero_24__22_  = \xz.mem_with_zero_24__22__sv2v_reg ;
  assign \xz.mem_with_zero_24__21_  = \xz.mem_with_zero_24__21__sv2v_reg ;
  assign \xz.mem_with_zero_24__20_  = \xz.mem_with_zero_24__20__sv2v_reg ;
  assign \xz.mem_with_zero_24__19_  = \xz.mem_with_zero_24__19__sv2v_reg ;
  assign \xz.mem_with_zero_24__18_  = \xz.mem_with_zero_24__18__sv2v_reg ;
  assign \xz.mem_with_zero_24__17_  = \xz.mem_with_zero_24__17__sv2v_reg ;
  assign \xz.mem_with_zero_24__16_  = \xz.mem_with_zero_24__16__sv2v_reg ;
  assign \xz.mem_with_zero_24__15_  = \xz.mem_with_zero_24__15__sv2v_reg ;
  assign \xz.mem_with_zero_24__14_  = \xz.mem_with_zero_24__14__sv2v_reg ;
  assign \xz.mem_with_zero_24__13_  = \xz.mem_with_zero_24__13__sv2v_reg ;
  assign \xz.mem_with_zero_24__12_  = \xz.mem_with_zero_24__12__sv2v_reg ;
  assign \xz.mem_with_zero_24__11_  = \xz.mem_with_zero_24__11__sv2v_reg ;
  assign \xz.mem_with_zero_24__10_  = \xz.mem_with_zero_24__10__sv2v_reg ;
  assign \xz.mem_with_zero_24__9_  = \xz.mem_with_zero_24__9__sv2v_reg ;
  assign \xz.mem_with_zero_24__8_  = \xz.mem_with_zero_24__8__sv2v_reg ;
  assign \xz.mem_with_zero_24__7_  = \xz.mem_with_zero_24__7__sv2v_reg ;
  assign \xz.mem_with_zero_24__6_  = \xz.mem_with_zero_24__6__sv2v_reg ;
  assign \xz.mem_with_zero_24__5_  = \xz.mem_with_zero_24__5__sv2v_reg ;
  assign \xz.mem_with_zero_24__4_  = \xz.mem_with_zero_24__4__sv2v_reg ;
  assign \xz.mem_with_zero_24__3_  = \xz.mem_with_zero_24__3__sv2v_reg ;
  assign \xz.mem_with_zero_24__2_  = \xz.mem_with_zero_24__2__sv2v_reg ;
  assign \xz.mem_with_zero_24__1_  = \xz.mem_with_zero_24__1__sv2v_reg ;
  assign \xz.mem_with_zero_24__0_  = \xz.mem_with_zero_24__0__sv2v_reg ;
  assign \xz.mem_with_zero_23__31_  = \xz.mem_with_zero_23__31__sv2v_reg ;
  assign \xz.mem_with_zero_23__30_  = \xz.mem_with_zero_23__30__sv2v_reg ;
  assign \xz.mem_with_zero_23__29_  = \xz.mem_with_zero_23__29__sv2v_reg ;
  assign \xz.mem_with_zero_23__28_  = \xz.mem_with_zero_23__28__sv2v_reg ;
  assign \xz.mem_with_zero_23__27_  = \xz.mem_with_zero_23__27__sv2v_reg ;
  assign \xz.mem_with_zero_23__26_  = \xz.mem_with_zero_23__26__sv2v_reg ;
  assign \xz.mem_with_zero_23__25_  = \xz.mem_with_zero_23__25__sv2v_reg ;
  assign \xz.mem_with_zero_23__24_  = \xz.mem_with_zero_23__24__sv2v_reg ;
  assign \xz.mem_with_zero_23__23_  = \xz.mem_with_zero_23__23__sv2v_reg ;
  assign \xz.mem_with_zero_23__22_  = \xz.mem_with_zero_23__22__sv2v_reg ;
  assign \xz.mem_with_zero_23__21_  = \xz.mem_with_zero_23__21__sv2v_reg ;
  assign \xz.mem_with_zero_23__20_  = \xz.mem_with_zero_23__20__sv2v_reg ;
  assign \xz.mem_with_zero_23__19_  = \xz.mem_with_zero_23__19__sv2v_reg ;
  assign \xz.mem_with_zero_23__18_  = \xz.mem_with_zero_23__18__sv2v_reg ;
  assign \xz.mem_with_zero_23__17_  = \xz.mem_with_zero_23__17__sv2v_reg ;
  assign \xz.mem_with_zero_23__16_  = \xz.mem_with_zero_23__16__sv2v_reg ;
  assign \xz.mem_with_zero_23__15_  = \xz.mem_with_zero_23__15__sv2v_reg ;
  assign \xz.mem_with_zero_23__14_  = \xz.mem_with_zero_23__14__sv2v_reg ;
  assign \xz.mem_with_zero_23__13_  = \xz.mem_with_zero_23__13__sv2v_reg ;
  assign \xz.mem_with_zero_23__12_  = \xz.mem_with_zero_23__12__sv2v_reg ;
  assign \xz.mem_with_zero_23__11_  = \xz.mem_with_zero_23__11__sv2v_reg ;
  assign \xz.mem_with_zero_23__10_  = \xz.mem_with_zero_23__10__sv2v_reg ;
  assign \xz.mem_with_zero_23__9_  = \xz.mem_with_zero_23__9__sv2v_reg ;
  assign \xz.mem_with_zero_23__8_  = \xz.mem_with_zero_23__8__sv2v_reg ;
  assign \xz.mem_with_zero_23__7_  = \xz.mem_with_zero_23__7__sv2v_reg ;
  assign \xz.mem_with_zero_23__6_  = \xz.mem_with_zero_23__6__sv2v_reg ;
  assign \xz.mem_with_zero_23__5_  = \xz.mem_with_zero_23__5__sv2v_reg ;
  assign \xz.mem_with_zero_23__4_  = \xz.mem_with_zero_23__4__sv2v_reg ;
  assign \xz.mem_with_zero_23__3_  = \xz.mem_with_zero_23__3__sv2v_reg ;
  assign \xz.mem_with_zero_23__2_  = \xz.mem_with_zero_23__2__sv2v_reg ;
  assign \xz.mem_with_zero_23__1_  = \xz.mem_with_zero_23__1__sv2v_reg ;
  assign \xz.mem_with_zero_23__0_  = \xz.mem_with_zero_23__0__sv2v_reg ;
  assign \xz.mem_with_zero_22__31_  = \xz.mem_with_zero_22__31__sv2v_reg ;
  assign \xz.mem_with_zero_22__30_  = \xz.mem_with_zero_22__30__sv2v_reg ;
  assign \xz.mem_with_zero_22__29_  = \xz.mem_with_zero_22__29__sv2v_reg ;
  assign \xz.mem_with_zero_22__28_  = \xz.mem_with_zero_22__28__sv2v_reg ;
  assign \xz.mem_with_zero_22__27_  = \xz.mem_with_zero_22__27__sv2v_reg ;
  assign \xz.mem_with_zero_22__26_  = \xz.mem_with_zero_22__26__sv2v_reg ;
  assign \xz.mem_with_zero_22__25_  = \xz.mem_with_zero_22__25__sv2v_reg ;
  assign \xz.mem_with_zero_22__24_  = \xz.mem_with_zero_22__24__sv2v_reg ;
  assign \xz.mem_with_zero_22__23_  = \xz.mem_with_zero_22__23__sv2v_reg ;
  assign \xz.mem_with_zero_22__22_  = \xz.mem_with_zero_22__22__sv2v_reg ;
  assign \xz.mem_with_zero_22__21_  = \xz.mem_with_zero_22__21__sv2v_reg ;
  assign \xz.mem_with_zero_22__20_  = \xz.mem_with_zero_22__20__sv2v_reg ;
  assign \xz.mem_with_zero_22__19_  = \xz.mem_with_zero_22__19__sv2v_reg ;
  assign \xz.mem_with_zero_22__18_  = \xz.mem_with_zero_22__18__sv2v_reg ;
  assign \xz.mem_with_zero_22__17_  = \xz.mem_with_zero_22__17__sv2v_reg ;
  assign \xz.mem_with_zero_22__16_  = \xz.mem_with_zero_22__16__sv2v_reg ;
  assign \xz.mem_with_zero_22__15_  = \xz.mem_with_zero_22__15__sv2v_reg ;
  assign \xz.mem_with_zero_22__14_  = \xz.mem_with_zero_22__14__sv2v_reg ;
  assign \xz.mem_with_zero_22__13_  = \xz.mem_with_zero_22__13__sv2v_reg ;
  assign \xz.mem_with_zero_22__12_  = \xz.mem_with_zero_22__12__sv2v_reg ;
  assign \xz.mem_with_zero_22__11_  = \xz.mem_with_zero_22__11__sv2v_reg ;
  assign \xz.mem_with_zero_22__10_  = \xz.mem_with_zero_22__10__sv2v_reg ;
  assign \xz.mem_with_zero_22__9_  = \xz.mem_with_zero_22__9__sv2v_reg ;
  assign \xz.mem_with_zero_22__8_  = \xz.mem_with_zero_22__8__sv2v_reg ;
  assign \xz.mem_with_zero_22__7_  = \xz.mem_with_zero_22__7__sv2v_reg ;
  assign \xz.mem_with_zero_22__6_  = \xz.mem_with_zero_22__6__sv2v_reg ;
  assign \xz.mem_with_zero_22__5_  = \xz.mem_with_zero_22__5__sv2v_reg ;
  assign \xz.mem_with_zero_22__4_  = \xz.mem_with_zero_22__4__sv2v_reg ;
  assign \xz.mem_with_zero_22__3_  = \xz.mem_with_zero_22__3__sv2v_reg ;
  assign \xz.mem_with_zero_22__2_  = \xz.mem_with_zero_22__2__sv2v_reg ;
  assign \xz.mem_with_zero_22__1_  = \xz.mem_with_zero_22__1__sv2v_reg ;
  assign \xz.mem_with_zero_22__0_  = \xz.mem_with_zero_22__0__sv2v_reg ;
  assign \xz.mem_with_zero_21__31_  = \xz.mem_with_zero_21__31__sv2v_reg ;
  assign \xz.mem_with_zero_21__30_  = \xz.mem_with_zero_21__30__sv2v_reg ;
  assign \xz.mem_with_zero_21__29_  = \xz.mem_with_zero_21__29__sv2v_reg ;
  assign \xz.mem_with_zero_21__28_  = \xz.mem_with_zero_21__28__sv2v_reg ;
  assign \xz.mem_with_zero_21__27_  = \xz.mem_with_zero_21__27__sv2v_reg ;
  assign \xz.mem_with_zero_21__26_  = \xz.mem_with_zero_21__26__sv2v_reg ;
  assign \xz.mem_with_zero_21__25_  = \xz.mem_with_zero_21__25__sv2v_reg ;
  assign \xz.mem_with_zero_21__24_  = \xz.mem_with_zero_21__24__sv2v_reg ;
  assign \xz.mem_with_zero_21__23_  = \xz.mem_with_zero_21__23__sv2v_reg ;
  assign \xz.mem_with_zero_21__22_  = \xz.mem_with_zero_21__22__sv2v_reg ;
  assign \xz.mem_with_zero_21__21_  = \xz.mem_with_zero_21__21__sv2v_reg ;
  assign \xz.mem_with_zero_21__20_  = \xz.mem_with_zero_21__20__sv2v_reg ;
  assign \xz.mem_with_zero_21__19_  = \xz.mem_with_zero_21__19__sv2v_reg ;
  assign \xz.mem_with_zero_21__18_  = \xz.mem_with_zero_21__18__sv2v_reg ;
  assign \xz.mem_with_zero_21__17_  = \xz.mem_with_zero_21__17__sv2v_reg ;
  assign \xz.mem_with_zero_21__16_  = \xz.mem_with_zero_21__16__sv2v_reg ;
  assign \xz.mem_with_zero_21__15_  = \xz.mem_with_zero_21__15__sv2v_reg ;
  assign \xz.mem_with_zero_21__14_  = \xz.mem_with_zero_21__14__sv2v_reg ;
  assign \xz.mem_with_zero_21__13_  = \xz.mem_with_zero_21__13__sv2v_reg ;
  assign \xz.mem_with_zero_21__12_  = \xz.mem_with_zero_21__12__sv2v_reg ;
  assign \xz.mem_with_zero_21__11_  = \xz.mem_with_zero_21__11__sv2v_reg ;
  assign \xz.mem_with_zero_21__10_  = \xz.mem_with_zero_21__10__sv2v_reg ;
  assign \xz.mem_with_zero_21__9_  = \xz.mem_with_zero_21__9__sv2v_reg ;
  assign \xz.mem_with_zero_21__8_  = \xz.mem_with_zero_21__8__sv2v_reg ;
  assign \xz.mem_with_zero_21__7_  = \xz.mem_with_zero_21__7__sv2v_reg ;
  assign \xz.mem_with_zero_21__6_  = \xz.mem_with_zero_21__6__sv2v_reg ;
  assign \xz.mem_with_zero_21__5_  = \xz.mem_with_zero_21__5__sv2v_reg ;
  assign \xz.mem_with_zero_21__4_  = \xz.mem_with_zero_21__4__sv2v_reg ;
  assign \xz.mem_with_zero_21__3_  = \xz.mem_with_zero_21__3__sv2v_reg ;
  assign \xz.mem_with_zero_21__2_  = \xz.mem_with_zero_21__2__sv2v_reg ;
  assign \xz.mem_with_zero_21__1_  = \xz.mem_with_zero_21__1__sv2v_reg ;
  assign \xz.mem_with_zero_21__0_  = \xz.mem_with_zero_21__0__sv2v_reg ;
  assign \xz.mem_with_zero_20__31_  = \xz.mem_with_zero_20__31__sv2v_reg ;
  assign \xz.mem_with_zero_20__30_  = \xz.mem_with_zero_20__30__sv2v_reg ;
  assign \xz.mem_with_zero_20__29_  = \xz.mem_with_zero_20__29__sv2v_reg ;
  assign \xz.mem_with_zero_20__28_  = \xz.mem_with_zero_20__28__sv2v_reg ;
  assign \xz.mem_with_zero_20__27_  = \xz.mem_with_zero_20__27__sv2v_reg ;
  assign \xz.mem_with_zero_20__26_  = \xz.mem_with_zero_20__26__sv2v_reg ;
  assign \xz.mem_with_zero_20__25_  = \xz.mem_with_zero_20__25__sv2v_reg ;
  assign \xz.mem_with_zero_20__24_  = \xz.mem_with_zero_20__24__sv2v_reg ;
  assign \xz.mem_with_zero_20__23_  = \xz.mem_with_zero_20__23__sv2v_reg ;
  assign \xz.mem_with_zero_20__22_  = \xz.mem_with_zero_20__22__sv2v_reg ;
  assign \xz.mem_with_zero_20__21_  = \xz.mem_with_zero_20__21__sv2v_reg ;
  assign \xz.mem_with_zero_20__20_  = \xz.mem_with_zero_20__20__sv2v_reg ;
  assign \xz.mem_with_zero_20__19_  = \xz.mem_with_zero_20__19__sv2v_reg ;
  assign \xz.mem_with_zero_20__18_  = \xz.mem_with_zero_20__18__sv2v_reg ;
  assign \xz.mem_with_zero_20__17_  = \xz.mem_with_zero_20__17__sv2v_reg ;
  assign \xz.mem_with_zero_20__16_  = \xz.mem_with_zero_20__16__sv2v_reg ;
  assign \xz.mem_with_zero_20__15_  = \xz.mem_with_zero_20__15__sv2v_reg ;
  assign \xz.mem_with_zero_20__14_  = \xz.mem_with_zero_20__14__sv2v_reg ;
  assign \xz.mem_with_zero_20__13_  = \xz.mem_with_zero_20__13__sv2v_reg ;
  assign \xz.mem_with_zero_20__12_  = \xz.mem_with_zero_20__12__sv2v_reg ;
  assign \xz.mem_with_zero_20__11_  = \xz.mem_with_zero_20__11__sv2v_reg ;
  assign \xz.mem_with_zero_20__10_  = \xz.mem_with_zero_20__10__sv2v_reg ;
  assign \xz.mem_with_zero_20__9_  = \xz.mem_with_zero_20__9__sv2v_reg ;
  assign \xz.mem_with_zero_20__8_  = \xz.mem_with_zero_20__8__sv2v_reg ;
  assign \xz.mem_with_zero_20__7_  = \xz.mem_with_zero_20__7__sv2v_reg ;
  assign \xz.mem_with_zero_20__6_  = \xz.mem_with_zero_20__6__sv2v_reg ;
  assign \xz.mem_with_zero_20__5_  = \xz.mem_with_zero_20__5__sv2v_reg ;
  assign \xz.mem_with_zero_20__4_  = \xz.mem_with_zero_20__4__sv2v_reg ;
  assign \xz.mem_with_zero_20__3_  = \xz.mem_with_zero_20__3__sv2v_reg ;
  assign \xz.mem_with_zero_20__2_  = \xz.mem_with_zero_20__2__sv2v_reg ;
  assign \xz.mem_with_zero_20__1_  = \xz.mem_with_zero_20__1__sv2v_reg ;
  assign \xz.mem_with_zero_20__0_  = \xz.mem_with_zero_20__0__sv2v_reg ;
  assign \xz.mem_with_zero_19__31_  = \xz.mem_with_zero_19__31__sv2v_reg ;
  assign \xz.mem_with_zero_19__30_  = \xz.mem_with_zero_19__30__sv2v_reg ;
  assign \xz.mem_with_zero_19__29_  = \xz.mem_with_zero_19__29__sv2v_reg ;
  assign \xz.mem_with_zero_19__28_  = \xz.mem_with_zero_19__28__sv2v_reg ;
  assign \xz.mem_with_zero_19__27_  = \xz.mem_with_zero_19__27__sv2v_reg ;
  assign \xz.mem_with_zero_19__26_  = \xz.mem_with_zero_19__26__sv2v_reg ;
  assign \xz.mem_with_zero_19__25_  = \xz.mem_with_zero_19__25__sv2v_reg ;
  assign \xz.mem_with_zero_19__24_  = \xz.mem_with_zero_19__24__sv2v_reg ;
  assign \xz.mem_with_zero_19__23_  = \xz.mem_with_zero_19__23__sv2v_reg ;
  assign \xz.mem_with_zero_19__22_  = \xz.mem_with_zero_19__22__sv2v_reg ;
  assign \xz.mem_with_zero_19__21_  = \xz.mem_with_zero_19__21__sv2v_reg ;
  assign \xz.mem_with_zero_19__20_  = \xz.mem_with_zero_19__20__sv2v_reg ;
  assign \xz.mem_with_zero_19__19_  = \xz.mem_with_zero_19__19__sv2v_reg ;
  assign \xz.mem_with_zero_19__18_  = \xz.mem_with_zero_19__18__sv2v_reg ;
  assign \xz.mem_with_zero_19__17_  = \xz.mem_with_zero_19__17__sv2v_reg ;
  assign \xz.mem_with_zero_19__16_  = \xz.mem_with_zero_19__16__sv2v_reg ;
  assign \xz.mem_with_zero_19__15_  = \xz.mem_with_zero_19__15__sv2v_reg ;
  assign \xz.mem_with_zero_19__14_  = \xz.mem_with_zero_19__14__sv2v_reg ;
  assign \xz.mem_with_zero_19__13_  = \xz.mem_with_zero_19__13__sv2v_reg ;
  assign \xz.mem_with_zero_19__12_  = \xz.mem_with_zero_19__12__sv2v_reg ;
  assign \xz.mem_with_zero_19__11_  = \xz.mem_with_zero_19__11__sv2v_reg ;
  assign \xz.mem_with_zero_19__10_  = \xz.mem_with_zero_19__10__sv2v_reg ;
  assign \xz.mem_with_zero_19__9_  = \xz.mem_with_zero_19__9__sv2v_reg ;
  assign \xz.mem_with_zero_19__8_  = \xz.mem_with_zero_19__8__sv2v_reg ;
  assign \xz.mem_with_zero_19__7_  = \xz.mem_with_zero_19__7__sv2v_reg ;
  assign \xz.mem_with_zero_19__6_  = \xz.mem_with_zero_19__6__sv2v_reg ;
  assign \xz.mem_with_zero_19__5_  = \xz.mem_with_zero_19__5__sv2v_reg ;
  assign \xz.mem_with_zero_19__4_  = \xz.mem_with_zero_19__4__sv2v_reg ;
  assign \xz.mem_with_zero_19__3_  = \xz.mem_with_zero_19__3__sv2v_reg ;
  assign \xz.mem_with_zero_19__2_  = \xz.mem_with_zero_19__2__sv2v_reg ;
  assign \xz.mem_with_zero_19__1_  = \xz.mem_with_zero_19__1__sv2v_reg ;
  assign \xz.mem_with_zero_19__0_  = \xz.mem_with_zero_19__0__sv2v_reg ;
  assign \xz.mem_with_zero_18__31_  = \xz.mem_with_zero_18__31__sv2v_reg ;
  assign \xz.mem_with_zero_18__30_  = \xz.mem_with_zero_18__30__sv2v_reg ;
  assign \xz.mem_with_zero_18__29_  = \xz.mem_with_zero_18__29__sv2v_reg ;
  assign \xz.mem_with_zero_18__28_  = \xz.mem_with_zero_18__28__sv2v_reg ;
  assign \xz.mem_with_zero_18__27_  = \xz.mem_with_zero_18__27__sv2v_reg ;
  assign \xz.mem_with_zero_18__26_  = \xz.mem_with_zero_18__26__sv2v_reg ;
  assign \xz.mem_with_zero_18__25_  = \xz.mem_with_zero_18__25__sv2v_reg ;
  assign \xz.mem_with_zero_18__24_  = \xz.mem_with_zero_18__24__sv2v_reg ;
  assign \xz.mem_with_zero_18__23_  = \xz.mem_with_zero_18__23__sv2v_reg ;
  assign \xz.mem_with_zero_18__22_  = \xz.mem_with_zero_18__22__sv2v_reg ;
  assign \xz.mem_with_zero_18__21_  = \xz.mem_with_zero_18__21__sv2v_reg ;
  assign \xz.mem_with_zero_18__20_  = \xz.mem_with_zero_18__20__sv2v_reg ;
  assign \xz.mem_with_zero_18__19_  = \xz.mem_with_zero_18__19__sv2v_reg ;
  assign \xz.mem_with_zero_18__18_  = \xz.mem_with_zero_18__18__sv2v_reg ;
  assign \xz.mem_with_zero_18__17_  = \xz.mem_with_zero_18__17__sv2v_reg ;
  assign \xz.mem_with_zero_18__16_  = \xz.mem_with_zero_18__16__sv2v_reg ;
  assign \xz.mem_with_zero_18__15_  = \xz.mem_with_zero_18__15__sv2v_reg ;
  assign \xz.mem_with_zero_18__14_  = \xz.mem_with_zero_18__14__sv2v_reg ;
  assign \xz.mem_with_zero_18__13_  = \xz.mem_with_zero_18__13__sv2v_reg ;
  assign \xz.mem_with_zero_18__12_  = \xz.mem_with_zero_18__12__sv2v_reg ;
  assign \xz.mem_with_zero_18__11_  = \xz.mem_with_zero_18__11__sv2v_reg ;
  assign \xz.mem_with_zero_18__10_  = \xz.mem_with_zero_18__10__sv2v_reg ;
  assign \xz.mem_with_zero_18__9_  = \xz.mem_with_zero_18__9__sv2v_reg ;
  assign \xz.mem_with_zero_18__8_  = \xz.mem_with_zero_18__8__sv2v_reg ;
  assign \xz.mem_with_zero_18__7_  = \xz.mem_with_zero_18__7__sv2v_reg ;
  assign \xz.mem_with_zero_18__6_  = \xz.mem_with_zero_18__6__sv2v_reg ;
  assign \xz.mem_with_zero_18__5_  = \xz.mem_with_zero_18__5__sv2v_reg ;
  assign \xz.mem_with_zero_18__4_  = \xz.mem_with_zero_18__4__sv2v_reg ;
  assign \xz.mem_with_zero_18__3_  = \xz.mem_with_zero_18__3__sv2v_reg ;
  assign \xz.mem_with_zero_18__2_  = \xz.mem_with_zero_18__2__sv2v_reg ;
  assign \xz.mem_with_zero_18__1_  = \xz.mem_with_zero_18__1__sv2v_reg ;
  assign \xz.mem_with_zero_18__0_  = \xz.mem_with_zero_18__0__sv2v_reg ;
  assign \xz.mem_with_zero_17__31_  = \xz.mem_with_zero_17__31__sv2v_reg ;
  assign \xz.mem_with_zero_17__30_  = \xz.mem_with_zero_17__30__sv2v_reg ;
  assign \xz.mem_with_zero_17__29_  = \xz.mem_with_zero_17__29__sv2v_reg ;
  assign \xz.mem_with_zero_17__28_  = \xz.mem_with_zero_17__28__sv2v_reg ;
  assign \xz.mem_with_zero_17__27_  = \xz.mem_with_zero_17__27__sv2v_reg ;
  assign \xz.mem_with_zero_17__26_  = \xz.mem_with_zero_17__26__sv2v_reg ;
  assign \xz.mem_with_zero_17__25_  = \xz.mem_with_zero_17__25__sv2v_reg ;
  assign \xz.mem_with_zero_17__24_  = \xz.mem_with_zero_17__24__sv2v_reg ;
  assign \xz.mem_with_zero_17__23_  = \xz.mem_with_zero_17__23__sv2v_reg ;
  assign \xz.mem_with_zero_17__22_  = \xz.mem_with_zero_17__22__sv2v_reg ;
  assign \xz.mem_with_zero_17__21_  = \xz.mem_with_zero_17__21__sv2v_reg ;
  assign \xz.mem_with_zero_17__20_  = \xz.mem_with_zero_17__20__sv2v_reg ;
  assign \xz.mem_with_zero_17__19_  = \xz.mem_with_zero_17__19__sv2v_reg ;
  assign \xz.mem_with_zero_17__18_  = \xz.mem_with_zero_17__18__sv2v_reg ;
  assign \xz.mem_with_zero_17__17_  = \xz.mem_with_zero_17__17__sv2v_reg ;
  assign \xz.mem_with_zero_17__16_  = \xz.mem_with_zero_17__16__sv2v_reg ;
  assign \xz.mem_with_zero_17__15_  = \xz.mem_with_zero_17__15__sv2v_reg ;
  assign \xz.mem_with_zero_17__14_  = \xz.mem_with_zero_17__14__sv2v_reg ;
  assign \xz.mem_with_zero_17__13_  = \xz.mem_with_zero_17__13__sv2v_reg ;
  assign \xz.mem_with_zero_17__12_  = \xz.mem_with_zero_17__12__sv2v_reg ;
  assign \xz.mem_with_zero_17__11_  = \xz.mem_with_zero_17__11__sv2v_reg ;
  assign \xz.mem_with_zero_17__10_  = \xz.mem_with_zero_17__10__sv2v_reg ;
  assign \xz.mem_with_zero_17__9_  = \xz.mem_with_zero_17__9__sv2v_reg ;
  assign \xz.mem_with_zero_17__8_  = \xz.mem_with_zero_17__8__sv2v_reg ;
  assign \xz.mem_with_zero_17__7_  = \xz.mem_with_zero_17__7__sv2v_reg ;
  assign \xz.mem_with_zero_17__6_  = \xz.mem_with_zero_17__6__sv2v_reg ;
  assign \xz.mem_with_zero_17__5_  = \xz.mem_with_zero_17__5__sv2v_reg ;
  assign \xz.mem_with_zero_17__4_  = \xz.mem_with_zero_17__4__sv2v_reg ;
  assign \xz.mem_with_zero_17__3_  = \xz.mem_with_zero_17__3__sv2v_reg ;
  assign \xz.mem_with_zero_17__2_  = \xz.mem_with_zero_17__2__sv2v_reg ;
  assign \xz.mem_with_zero_17__1_  = \xz.mem_with_zero_17__1__sv2v_reg ;
  assign \xz.mem_with_zero_17__0_  = \xz.mem_with_zero_17__0__sv2v_reg ;
  assign \xz.mem_with_zero_16__31_  = \xz.mem_with_zero_16__31__sv2v_reg ;
  assign \xz.mem_with_zero_16__30_  = \xz.mem_with_zero_16__30__sv2v_reg ;
  assign \xz.mem_with_zero_16__29_  = \xz.mem_with_zero_16__29__sv2v_reg ;
  assign \xz.mem_with_zero_16__28_  = \xz.mem_with_zero_16__28__sv2v_reg ;
  assign \xz.mem_with_zero_16__27_  = \xz.mem_with_zero_16__27__sv2v_reg ;
  assign \xz.mem_with_zero_16__26_  = \xz.mem_with_zero_16__26__sv2v_reg ;
  assign \xz.mem_with_zero_16__25_  = \xz.mem_with_zero_16__25__sv2v_reg ;
  assign \xz.mem_with_zero_16__24_  = \xz.mem_with_zero_16__24__sv2v_reg ;
  assign \xz.mem_with_zero_16__23_  = \xz.mem_with_zero_16__23__sv2v_reg ;
  assign \xz.mem_with_zero_16__22_  = \xz.mem_with_zero_16__22__sv2v_reg ;
  assign \xz.mem_with_zero_16__21_  = \xz.mem_with_zero_16__21__sv2v_reg ;
  assign \xz.mem_with_zero_16__20_  = \xz.mem_with_zero_16__20__sv2v_reg ;
  assign \xz.mem_with_zero_16__19_  = \xz.mem_with_zero_16__19__sv2v_reg ;
  assign \xz.mem_with_zero_16__18_  = \xz.mem_with_zero_16__18__sv2v_reg ;
  assign \xz.mem_with_zero_16__17_  = \xz.mem_with_zero_16__17__sv2v_reg ;
  assign \xz.mem_with_zero_16__16_  = \xz.mem_with_zero_16__16__sv2v_reg ;
  assign \xz.mem_with_zero_16__15_  = \xz.mem_with_zero_16__15__sv2v_reg ;
  assign \xz.mem_with_zero_16__14_  = \xz.mem_with_zero_16__14__sv2v_reg ;
  assign \xz.mem_with_zero_16__13_  = \xz.mem_with_zero_16__13__sv2v_reg ;
  assign \xz.mem_with_zero_16__12_  = \xz.mem_with_zero_16__12__sv2v_reg ;
  assign \xz.mem_with_zero_16__11_  = \xz.mem_with_zero_16__11__sv2v_reg ;
  assign \xz.mem_with_zero_16__10_  = \xz.mem_with_zero_16__10__sv2v_reg ;
  assign \xz.mem_with_zero_16__9_  = \xz.mem_with_zero_16__9__sv2v_reg ;
  assign \xz.mem_with_zero_16__8_  = \xz.mem_with_zero_16__8__sv2v_reg ;
  assign \xz.mem_with_zero_16__7_  = \xz.mem_with_zero_16__7__sv2v_reg ;
  assign \xz.mem_with_zero_16__6_  = \xz.mem_with_zero_16__6__sv2v_reg ;
  assign \xz.mem_with_zero_16__5_  = \xz.mem_with_zero_16__5__sv2v_reg ;
  assign \xz.mem_with_zero_16__4_  = \xz.mem_with_zero_16__4__sv2v_reg ;
  assign \xz.mem_with_zero_16__3_  = \xz.mem_with_zero_16__3__sv2v_reg ;
  assign \xz.mem_with_zero_16__2_  = \xz.mem_with_zero_16__2__sv2v_reg ;
  assign \xz.mem_with_zero_16__1_  = \xz.mem_with_zero_16__1__sv2v_reg ;
  assign \xz.mem_with_zero_16__0_  = \xz.mem_with_zero_16__0__sv2v_reg ;
  assign \xz.mem_with_zero_15__31_  = \xz.mem_with_zero_15__31__sv2v_reg ;
  assign \xz.mem_with_zero_15__30_  = \xz.mem_with_zero_15__30__sv2v_reg ;
  assign \xz.mem_with_zero_15__29_  = \xz.mem_with_zero_15__29__sv2v_reg ;
  assign \xz.mem_with_zero_15__28_  = \xz.mem_with_zero_15__28__sv2v_reg ;
  assign \xz.mem_with_zero_15__27_  = \xz.mem_with_zero_15__27__sv2v_reg ;
  assign \xz.mem_with_zero_15__26_  = \xz.mem_with_zero_15__26__sv2v_reg ;
  assign \xz.mem_with_zero_15__25_  = \xz.mem_with_zero_15__25__sv2v_reg ;
  assign \xz.mem_with_zero_15__24_  = \xz.mem_with_zero_15__24__sv2v_reg ;
  assign \xz.mem_with_zero_15__23_  = \xz.mem_with_zero_15__23__sv2v_reg ;
  assign \xz.mem_with_zero_15__22_  = \xz.mem_with_zero_15__22__sv2v_reg ;
  assign \xz.mem_with_zero_15__21_  = \xz.mem_with_zero_15__21__sv2v_reg ;
  assign \xz.mem_with_zero_15__20_  = \xz.mem_with_zero_15__20__sv2v_reg ;
  assign \xz.mem_with_zero_15__19_  = \xz.mem_with_zero_15__19__sv2v_reg ;
  assign \xz.mem_with_zero_15__18_  = \xz.mem_with_zero_15__18__sv2v_reg ;
  assign \xz.mem_with_zero_15__17_  = \xz.mem_with_zero_15__17__sv2v_reg ;
  assign \xz.mem_with_zero_15__16_  = \xz.mem_with_zero_15__16__sv2v_reg ;
  assign \xz.mem_with_zero_15__15_  = \xz.mem_with_zero_15__15__sv2v_reg ;
  assign \xz.mem_with_zero_15__14_  = \xz.mem_with_zero_15__14__sv2v_reg ;
  assign \xz.mem_with_zero_15__13_  = \xz.mem_with_zero_15__13__sv2v_reg ;
  assign \xz.mem_with_zero_15__12_  = \xz.mem_with_zero_15__12__sv2v_reg ;
  assign \xz.mem_with_zero_15__11_  = \xz.mem_with_zero_15__11__sv2v_reg ;
  assign \xz.mem_with_zero_15__10_  = \xz.mem_with_zero_15__10__sv2v_reg ;
  assign \xz.mem_with_zero_15__9_  = \xz.mem_with_zero_15__9__sv2v_reg ;
  assign \xz.mem_with_zero_15__8_  = \xz.mem_with_zero_15__8__sv2v_reg ;
  assign \xz.mem_with_zero_15__7_  = \xz.mem_with_zero_15__7__sv2v_reg ;
  assign \xz.mem_with_zero_15__6_  = \xz.mem_with_zero_15__6__sv2v_reg ;
  assign \xz.mem_with_zero_15__5_  = \xz.mem_with_zero_15__5__sv2v_reg ;
  assign \xz.mem_with_zero_15__4_  = \xz.mem_with_zero_15__4__sv2v_reg ;
  assign \xz.mem_with_zero_15__3_  = \xz.mem_with_zero_15__3__sv2v_reg ;
  assign \xz.mem_with_zero_15__2_  = \xz.mem_with_zero_15__2__sv2v_reg ;
  assign \xz.mem_with_zero_15__1_  = \xz.mem_with_zero_15__1__sv2v_reg ;
  assign \xz.mem_with_zero_15__0_  = \xz.mem_with_zero_15__0__sv2v_reg ;
  assign \xz.mem_with_zero_14__31_  = \xz.mem_with_zero_14__31__sv2v_reg ;
  assign \xz.mem_with_zero_14__30_  = \xz.mem_with_zero_14__30__sv2v_reg ;
  assign \xz.mem_with_zero_14__29_  = \xz.mem_with_zero_14__29__sv2v_reg ;
  assign \xz.mem_with_zero_14__28_  = \xz.mem_with_zero_14__28__sv2v_reg ;
  assign \xz.mem_with_zero_14__27_  = \xz.mem_with_zero_14__27__sv2v_reg ;
  assign \xz.mem_with_zero_14__26_  = \xz.mem_with_zero_14__26__sv2v_reg ;
  assign \xz.mem_with_zero_14__25_  = \xz.mem_with_zero_14__25__sv2v_reg ;
  assign \xz.mem_with_zero_14__24_  = \xz.mem_with_zero_14__24__sv2v_reg ;
  assign \xz.mem_with_zero_14__23_  = \xz.mem_with_zero_14__23__sv2v_reg ;
  assign \xz.mem_with_zero_14__22_  = \xz.mem_with_zero_14__22__sv2v_reg ;
  assign \xz.mem_with_zero_14__21_  = \xz.mem_with_zero_14__21__sv2v_reg ;
  assign \xz.mem_with_zero_14__20_  = \xz.mem_with_zero_14__20__sv2v_reg ;
  assign \xz.mem_with_zero_14__19_  = \xz.mem_with_zero_14__19__sv2v_reg ;
  assign \xz.mem_with_zero_14__18_  = \xz.mem_with_zero_14__18__sv2v_reg ;
  assign \xz.mem_with_zero_14__17_  = \xz.mem_with_zero_14__17__sv2v_reg ;
  assign \xz.mem_with_zero_14__16_  = \xz.mem_with_zero_14__16__sv2v_reg ;
  assign \xz.mem_with_zero_14__15_  = \xz.mem_with_zero_14__15__sv2v_reg ;
  assign \xz.mem_with_zero_14__14_  = \xz.mem_with_zero_14__14__sv2v_reg ;
  assign \xz.mem_with_zero_14__13_  = \xz.mem_with_zero_14__13__sv2v_reg ;
  assign \xz.mem_with_zero_14__12_  = \xz.mem_with_zero_14__12__sv2v_reg ;
  assign \xz.mem_with_zero_14__11_  = \xz.mem_with_zero_14__11__sv2v_reg ;
  assign \xz.mem_with_zero_14__10_  = \xz.mem_with_zero_14__10__sv2v_reg ;
  assign \xz.mem_with_zero_14__9_  = \xz.mem_with_zero_14__9__sv2v_reg ;
  assign \xz.mem_with_zero_14__8_  = \xz.mem_with_zero_14__8__sv2v_reg ;
  assign \xz.mem_with_zero_14__7_  = \xz.mem_with_zero_14__7__sv2v_reg ;
  assign \xz.mem_with_zero_14__6_  = \xz.mem_with_zero_14__6__sv2v_reg ;
  assign \xz.mem_with_zero_14__5_  = \xz.mem_with_zero_14__5__sv2v_reg ;
  assign \xz.mem_with_zero_14__4_  = \xz.mem_with_zero_14__4__sv2v_reg ;
  assign \xz.mem_with_zero_14__3_  = \xz.mem_with_zero_14__3__sv2v_reg ;
  assign \xz.mem_with_zero_14__2_  = \xz.mem_with_zero_14__2__sv2v_reg ;
  assign \xz.mem_with_zero_14__1_  = \xz.mem_with_zero_14__1__sv2v_reg ;
  assign \xz.mem_with_zero_14__0_  = \xz.mem_with_zero_14__0__sv2v_reg ;
  assign \xz.mem_with_zero_13__31_  = \xz.mem_with_zero_13__31__sv2v_reg ;
  assign \xz.mem_with_zero_13__30_  = \xz.mem_with_zero_13__30__sv2v_reg ;
  assign \xz.mem_with_zero_13__29_  = \xz.mem_with_zero_13__29__sv2v_reg ;
  assign \xz.mem_with_zero_13__28_  = \xz.mem_with_zero_13__28__sv2v_reg ;
  assign \xz.mem_with_zero_13__27_  = \xz.mem_with_zero_13__27__sv2v_reg ;
  assign \xz.mem_with_zero_13__26_  = \xz.mem_with_zero_13__26__sv2v_reg ;
  assign \xz.mem_with_zero_13__25_  = \xz.mem_with_zero_13__25__sv2v_reg ;
  assign \xz.mem_with_zero_13__24_  = \xz.mem_with_zero_13__24__sv2v_reg ;
  assign \xz.mem_with_zero_13__23_  = \xz.mem_with_zero_13__23__sv2v_reg ;
  assign \xz.mem_with_zero_13__22_  = \xz.mem_with_zero_13__22__sv2v_reg ;
  assign \xz.mem_with_zero_13__21_  = \xz.mem_with_zero_13__21__sv2v_reg ;
  assign \xz.mem_with_zero_13__20_  = \xz.mem_with_zero_13__20__sv2v_reg ;
  assign \xz.mem_with_zero_13__19_  = \xz.mem_with_zero_13__19__sv2v_reg ;
  assign \xz.mem_with_zero_13__18_  = \xz.mem_with_zero_13__18__sv2v_reg ;
  assign \xz.mem_with_zero_13__17_  = \xz.mem_with_zero_13__17__sv2v_reg ;
  assign \xz.mem_with_zero_13__16_  = \xz.mem_with_zero_13__16__sv2v_reg ;
  assign \xz.mem_with_zero_13__15_  = \xz.mem_with_zero_13__15__sv2v_reg ;
  assign \xz.mem_with_zero_13__14_  = \xz.mem_with_zero_13__14__sv2v_reg ;
  assign \xz.mem_with_zero_13__13_  = \xz.mem_with_zero_13__13__sv2v_reg ;
  assign \xz.mem_with_zero_13__12_  = \xz.mem_with_zero_13__12__sv2v_reg ;
  assign \xz.mem_with_zero_13__11_  = \xz.mem_with_zero_13__11__sv2v_reg ;
  assign \xz.mem_with_zero_13__10_  = \xz.mem_with_zero_13__10__sv2v_reg ;
  assign \xz.mem_with_zero_13__9_  = \xz.mem_with_zero_13__9__sv2v_reg ;
  assign \xz.mem_with_zero_13__8_  = \xz.mem_with_zero_13__8__sv2v_reg ;
  assign \xz.mem_with_zero_13__7_  = \xz.mem_with_zero_13__7__sv2v_reg ;
  assign \xz.mem_with_zero_13__6_  = \xz.mem_with_zero_13__6__sv2v_reg ;
  assign \xz.mem_with_zero_13__5_  = \xz.mem_with_zero_13__5__sv2v_reg ;
  assign \xz.mem_with_zero_13__4_  = \xz.mem_with_zero_13__4__sv2v_reg ;
  assign \xz.mem_with_zero_13__3_  = \xz.mem_with_zero_13__3__sv2v_reg ;
  assign \xz.mem_with_zero_13__2_  = \xz.mem_with_zero_13__2__sv2v_reg ;
  assign \xz.mem_with_zero_13__1_  = \xz.mem_with_zero_13__1__sv2v_reg ;
  assign \xz.mem_with_zero_13__0_  = \xz.mem_with_zero_13__0__sv2v_reg ;
  assign \xz.mem_with_zero_12__31_  = \xz.mem_with_zero_12__31__sv2v_reg ;
  assign \xz.mem_with_zero_12__30_  = \xz.mem_with_zero_12__30__sv2v_reg ;
  assign \xz.mem_with_zero_12__29_  = \xz.mem_with_zero_12__29__sv2v_reg ;
  assign \xz.mem_with_zero_12__28_  = \xz.mem_with_zero_12__28__sv2v_reg ;
  assign \xz.mem_with_zero_12__27_  = \xz.mem_with_zero_12__27__sv2v_reg ;
  assign \xz.mem_with_zero_12__26_  = \xz.mem_with_zero_12__26__sv2v_reg ;
  assign \xz.mem_with_zero_12__25_  = \xz.mem_with_zero_12__25__sv2v_reg ;
  assign \xz.mem_with_zero_12__24_  = \xz.mem_with_zero_12__24__sv2v_reg ;
  assign \xz.mem_with_zero_12__23_  = \xz.mem_with_zero_12__23__sv2v_reg ;
  assign \xz.mem_with_zero_12__22_  = \xz.mem_with_zero_12__22__sv2v_reg ;
  assign \xz.mem_with_zero_12__21_  = \xz.mem_with_zero_12__21__sv2v_reg ;
  assign \xz.mem_with_zero_12__20_  = \xz.mem_with_zero_12__20__sv2v_reg ;
  assign \xz.mem_with_zero_12__19_  = \xz.mem_with_zero_12__19__sv2v_reg ;
  assign \xz.mem_with_zero_12__18_  = \xz.mem_with_zero_12__18__sv2v_reg ;
  assign \xz.mem_with_zero_12__17_  = \xz.mem_with_zero_12__17__sv2v_reg ;
  assign \xz.mem_with_zero_12__16_  = \xz.mem_with_zero_12__16__sv2v_reg ;
  assign \xz.mem_with_zero_12__15_  = \xz.mem_with_zero_12__15__sv2v_reg ;
  assign \xz.mem_with_zero_12__14_  = \xz.mem_with_zero_12__14__sv2v_reg ;
  assign \xz.mem_with_zero_12__13_  = \xz.mem_with_zero_12__13__sv2v_reg ;
  assign \xz.mem_with_zero_12__12_  = \xz.mem_with_zero_12__12__sv2v_reg ;
  assign \xz.mem_with_zero_12__11_  = \xz.mem_with_zero_12__11__sv2v_reg ;
  assign \xz.mem_with_zero_12__10_  = \xz.mem_with_zero_12__10__sv2v_reg ;
  assign \xz.mem_with_zero_12__9_  = \xz.mem_with_zero_12__9__sv2v_reg ;
  assign \xz.mem_with_zero_12__8_  = \xz.mem_with_zero_12__8__sv2v_reg ;
  assign \xz.mem_with_zero_12__7_  = \xz.mem_with_zero_12__7__sv2v_reg ;
  assign \xz.mem_with_zero_12__6_  = \xz.mem_with_zero_12__6__sv2v_reg ;
  assign \xz.mem_with_zero_12__5_  = \xz.mem_with_zero_12__5__sv2v_reg ;
  assign \xz.mem_with_zero_12__4_  = \xz.mem_with_zero_12__4__sv2v_reg ;
  assign \xz.mem_with_zero_12__3_  = \xz.mem_with_zero_12__3__sv2v_reg ;
  assign \xz.mem_with_zero_12__2_  = \xz.mem_with_zero_12__2__sv2v_reg ;
  assign \xz.mem_with_zero_12__1_  = \xz.mem_with_zero_12__1__sv2v_reg ;
  assign \xz.mem_with_zero_12__0_  = \xz.mem_with_zero_12__0__sv2v_reg ;
  assign \xz.mem_with_zero_11__31_  = \xz.mem_with_zero_11__31__sv2v_reg ;
  assign \xz.mem_with_zero_11__30_  = \xz.mem_with_zero_11__30__sv2v_reg ;
  assign \xz.mem_with_zero_11__29_  = \xz.mem_with_zero_11__29__sv2v_reg ;
  assign \xz.mem_with_zero_11__28_  = \xz.mem_with_zero_11__28__sv2v_reg ;
  assign \xz.mem_with_zero_11__27_  = \xz.mem_with_zero_11__27__sv2v_reg ;
  assign \xz.mem_with_zero_11__26_  = \xz.mem_with_zero_11__26__sv2v_reg ;
  assign \xz.mem_with_zero_11__25_  = \xz.mem_with_zero_11__25__sv2v_reg ;
  assign \xz.mem_with_zero_11__24_  = \xz.mem_with_zero_11__24__sv2v_reg ;
  assign \xz.mem_with_zero_11__23_  = \xz.mem_with_zero_11__23__sv2v_reg ;
  assign \xz.mem_with_zero_11__22_  = \xz.mem_with_zero_11__22__sv2v_reg ;
  assign \xz.mem_with_zero_11__21_  = \xz.mem_with_zero_11__21__sv2v_reg ;
  assign \xz.mem_with_zero_11__20_  = \xz.mem_with_zero_11__20__sv2v_reg ;
  assign \xz.mem_with_zero_11__19_  = \xz.mem_with_zero_11__19__sv2v_reg ;
  assign \xz.mem_with_zero_11__18_  = \xz.mem_with_zero_11__18__sv2v_reg ;
  assign \xz.mem_with_zero_11__17_  = \xz.mem_with_zero_11__17__sv2v_reg ;
  assign \xz.mem_with_zero_11__16_  = \xz.mem_with_zero_11__16__sv2v_reg ;
  assign \xz.mem_with_zero_11__15_  = \xz.mem_with_zero_11__15__sv2v_reg ;
  assign \xz.mem_with_zero_11__14_  = \xz.mem_with_zero_11__14__sv2v_reg ;
  assign \xz.mem_with_zero_11__13_  = \xz.mem_with_zero_11__13__sv2v_reg ;
  assign \xz.mem_with_zero_11__12_  = \xz.mem_with_zero_11__12__sv2v_reg ;
  assign \xz.mem_with_zero_11__11_  = \xz.mem_with_zero_11__11__sv2v_reg ;
  assign \xz.mem_with_zero_11__10_  = \xz.mem_with_zero_11__10__sv2v_reg ;
  assign \xz.mem_with_zero_11__9_  = \xz.mem_with_zero_11__9__sv2v_reg ;
  assign \xz.mem_with_zero_11__8_  = \xz.mem_with_zero_11__8__sv2v_reg ;
  assign \xz.mem_with_zero_11__7_  = \xz.mem_with_zero_11__7__sv2v_reg ;
  assign \xz.mem_with_zero_11__6_  = \xz.mem_with_zero_11__6__sv2v_reg ;
  assign \xz.mem_with_zero_11__5_  = \xz.mem_with_zero_11__5__sv2v_reg ;
  assign \xz.mem_with_zero_11__4_  = \xz.mem_with_zero_11__4__sv2v_reg ;
  assign \xz.mem_with_zero_11__3_  = \xz.mem_with_zero_11__3__sv2v_reg ;
  assign \xz.mem_with_zero_11__2_  = \xz.mem_with_zero_11__2__sv2v_reg ;
  assign \xz.mem_with_zero_11__1_  = \xz.mem_with_zero_11__1__sv2v_reg ;
  assign \xz.mem_with_zero_11__0_  = \xz.mem_with_zero_11__0__sv2v_reg ;
  assign \xz.mem_with_zero_10__31_  = \xz.mem_with_zero_10__31__sv2v_reg ;
  assign \xz.mem_with_zero_10__30_  = \xz.mem_with_zero_10__30__sv2v_reg ;
  assign \xz.mem_with_zero_10__29_  = \xz.mem_with_zero_10__29__sv2v_reg ;
  assign \xz.mem_with_zero_10__28_  = \xz.mem_with_zero_10__28__sv2v_reg ;
  assign \xz.mem_with_zero_10__27_  = \xz.mem_with_zero_10__27__sv2v_reg ;
  assign \xz.mem_with_zero_10__26_  = \xz.mem_with_zero_10__26__sv2v_reg ;
  assign \xz.mem_with_zero_10__25_  = \xz.mem_with_zero_10__25__sv2v_reg ;
  assign \xz.mem_with_zero_10__24_  = \xz.mem_with_zero_10__24__sv2v_reg ;
  assign \xz.mem_with_zero_10__23_  = \xz.mem_with_zero_10__23__sv2v_reg ;
  assign \xz.mem_with_zero_10__22_  = \xz.mem_with_zero_10__22__sv2v_reg ;
  assign \xz.mem_with_zero_10__21_  = \xz.mem_with_zero_10__21__sv2v_reg ;
  assign \xz.mem_with_zero_10__20_  = \xz.mem_with_zero_10__20__sv2v_reg ;
  assign \xz.mem_with_zero_10__19_  = \xz.mem_with_zero_10__19__sv2v_reg ;
  assign \xz.mem_with_zero_10__18_  = \xz.mem_with_zero_10__18__sv2v_reg ;
  assign \xz.mem_with_zero_10__17_  = \xz.mem_with_zero_10__17__sv2v_reg ;
  assign \xz.mem_with_zero_10__16_  = \xz.mem_with_zero_10__16__sv2v_reg ;
  assign \xz.mem_with_zero_10__15_  = \xz.mem_with_zero_10__15__sv2v_reg ;
  assign \xz.mem_with_zero_10__14_  = \xz.mem_with_zero_10__14__sv2v_reg ;
  assign \xz.mem_with_zero_10__13_  = \xz.mem_with_zero_10__13__sv2v_reg ;
  assign \xz.mem_with_zero_10__12_  = \xz.mem_with_zero_10__12__sv2v_reg ;
  assign \xz.mem_with_zero_10__11_  = \xz.mem_with_zero_10__11__sv2v_reg ;
  assign \xz.mem_with_zero_10__10_  = \xz.mem_with_zero_10__10__sv2v_reg ;
  assign \xz.mem_with_zero_10__9_  = \xz.mem_with_zero_10__9__sv2v_reg ;
  assign \xz.mem_with_zero_10__8_  = \xz.mem_with_zero_10__8__sv2v_reg ;
  assign \xz.mem_with_zero_10__7_  = \xz.mem_with_zero_10__7__sv2v_reg ;
  assign \xz.mem_with_zero_10__6_  = \xz.mem_with_zero_10__6__sv2v_reg ;
  assign \xz.mem_with_zero_10__5_  = \xz.mem_with_zero_10__5__sv2v_reg ;
  assign \xz.mem_with_zero_10__4_  = \xz.mem_with_zero_10__4__sv2v_reg ;
  assign \xz.mem_with_zero_10__3_  = \xz.mem_with_zero_10__3__sv2v_reg ;
  assign \xz.mem_with_zero_10__2_  = \xz.mem_with_zero_10__2__sv2v_reg ;
  assign \xz.mem_with_zero_10__1_  = \xz.mem_with_zero_10__1__sv2v_reg ;
  assign \xz.mem_with_zero_10__0_  = \xz.mem_with_zero_10__0__sv2v_reg ;
  assign \xz.mem_with_zero_9__31_  = \xz.mem_with_zero_9__31__sv2v_reg ;
  assign \xz.mem_with_zero_9__30_  = \xz.mem_with_zero_9__30__sv2v_reg ;
  assign \xz.mem_with_zero_9__29_  = \xz.mem_with_zero_9__29__sv2v_reg ;
  assign \xz.mem_with_zero_9__28_  = \xz.mem_with_zero_9__28__sv2v_reg ;
  assign \xz.mem_with_zero_9__27_  = \xz.mem_with_zero_9__27__sv2v_reg ;
  assign \xz.mem_with_zero_9__26_  = \xz.mem_with_zero_9__26__sv2v_reg ;
  assign \xz.mem_with_zero_9__25_  = \xz.mem_with_zero_9__25__sv2v_reg ;
  assign \xz.mem_with_zero_9__24_  = \xz.mem_with_zero_9__24__sv2v_reg ;
  assign \xz.mem_with_zero_9__23_  = \xz.mem_with_zero_9__23__sv2v_reg ;
  assign \xz.mem_with_zero_9__22_  = \xz.mem_with_zero_9__22__sv2v_reg ;
  assign \xz.mem_with_zero_9__21_  = \xz.mem_with_zero_9__21__sv2v_reg ;
  assign \xz.mem_with_zero_9__20_  = \xz.mem_with_zero_9__20__sv2v_reg ;
  assign \xz.mem_with_zero_9__19_  = \xz.mem_with_zero_9__19__sv2v_reg ;
  assign \xz.mem_with_zero_9__18_  = \xz.mem_with_zero_9__18__sv2v_reg ;
  assign \xz.mem_with_zero_9__17_  = \xz.mem_with_zero_9__17__sv2v_reg ;
  assign \xz.mem_with_zero_9__16_  = \xz.mem_with_zero_9__16__sv2v_reg ;
  assign \xz.mem_with_zero_9__15_  = \xz.mem_with_zero_9__15__sv2v_reg ;
  assign \xz.mem_with_zero_9__14_  = \xz.mem_with_zero_9__14__sv2v_reg ;
  assign \xz.mem_with_zero_9__13_  = \xz.mem_with_zero_9__13__sv2v_reg ;
  assign \xz.mem_with_zero_9__12_  = \xz.mem_with_zero_9__12__sv2v_reg ;
  assign \xz.mem_with_zero_9__11_  = \xz.mem_with_zero_9__11__sv2v_reg ;
  assign \xz.mem_with_zero_9__10_  = \xz.mem_with_zero_9__10__sv2v_reg ;
  assign \xz.mem_with_zero_9__9_  = \xz.mem_with_zero_9__9__sv2v_reg ;
  assign \xz.mem_with_zero_9__8_  = \xz.mem_with_zero_9__8__sv2v_reg ;
  assign \xz.mem_with_zero_9__7_  = \xz.mem_with_zero_9__7__sv2v_reg ;
  assign \xz.mem_with_zero_9__6_  = \xz.mem_with_zero_9__6__sv2v_reg ;
  assign \xz.mem_with_zero_9__5_  = \xz.mem_with_zero_9__5__sv2v_reg ;
  assign \xz.mem_with_zero_9__4_  = \xz.mem_with_zero_9__4__sv2v_reg ;
  assign \xz.mem_with_zero_9__3_  = \xz.mem_with_zero_9__3__sv2v_reg ;
  assign \xz.mem_with_zero_9__2_  = \xz.mem_with_zero_9__2__sv2v_reg ;
  assign \xz.mem_with_zero_9__1_  = \xz.mem_with_zero_9__1__sv2v_reg ;
  assign \xz.mem_with_zero_9__0_  = \xz.mem_with_zero_9__0__sv2v_reg ;
  assign \xz.mem_with_zero_8__31_  = \xz.mem_with_zero_8__31__sv2v_reg ;
  assign \xz.mem_with_zero_8__30_  = \xz.mem_with_zero_8__30__sv2v_reg ;
  assign \xz.mem_with_zero_8__29_  = \xz.mem_with_zero_8__29__sv2v_reg ;
  assign \xz.mem_with_zero_8__28_  = \xz.mem_with_zero_8__28__sv2v_reg ;
  assign \xz.mem_with_zero_8__27_  = \xz.mem_with_zero_8__27__sv2v_reg ;
  assign \xz.mem_with_zero_8__26_  = \xz.mem_with_zero_8__26__sv2v_reg ;
  assign \xz.mem_with_zero_8__25_  = \xz.mem_with_zero_8__25__sv2v_reg ;
  assign \xz.mem_with_zero_8__24_  = \xz.mem_with_zero_8__24__sv2v_reg ;
  assign \xz.mem_with_zero_8__23_  = \xz.mem_with_zero_8__23__sv2v_reg ;
  assign \xz.mem_with_zero_8__22_  = \xz.mem_with_zero_8__22__sv2v_reg ;
  assign \xz.mem_with_zero_8__21_  = \xz.mem_with_zero_8__21__sv2v_reg ;
  assign \xz.mem_with_zero_8__20_  = \xz.mem_with_zero_8__20__sv2v_reg ;
  assign \xz.mem_with_zero_8__19_  = \xz.mem_with_zero_8__19__sv2v_reg ;
  assign \xz.mem_with_zero_8__18_  = \xz.mem_with_zero_8__18__sv2v_reg ;
  assign \xz.mem_with_zero_8__17_  = \xz.mem_with_zero_8__17__sv2v_reg ;
  assign \xz.mem_with_zero_8__16_  = \xz.mem_with_zero_8__16__sv2v_reg ;
  assign \xz.mem_with_zero_8__15_  = \xz.mem_with_zero_8__15__sv2v_reg ;
  assign \xz.mem_with_zero_8__14_  = \xz.mem_with_zero_8__14__sv2v_reg ;
  assign \xz.mem_with_zero_8__13_  = \xz.mem_with_zero_8__13__sv2v_reg ;
  assign \xz.mem_with_zero_8__12_  = \xz.mem_with_zero_8__12__sv2v_reg ;
  assign \xz.mem_with_zero_8__11_  = \xz.mem_with_zero_8__11__sv2v_reg ;
  assign \xz.mem_with_zero_8__10_  = \xz.mem_with_zero_8__10__sv2v_reg ;
  assign \xz.mem_with_zero_8__9_  = \xz.mem_with_zero_8__9__sv2v_reg ;
  assign \xz.mem_with_zero_8__8_  = \xz.mem_with_zero_8__8__sv2v_reg ;
  assign \xz.mem_with_zero_8__7_  = \xz.mem_with_zero_8__7__sv2v_reg ;
  assign \xz.mem_with_zero_8__6_  = \xz.mem_with_zero_8__6__sv2v_reg ;
  assign \xz.mem_with_zero_8__5_  = \xz.mem_with_zero_8__5__sv2v_reg ;
  assign \xz.mem_with_zero_8__4_  = \xz.mem_with_zero_8__4__sv2v_reg ;
  assign \xz.mem_with_zero_8__3_  = \xz.mem_with_zero_8__3__sv2v_reg ;
  assign \xz.mem_with_zero_8__2_  = \xz.mem_with_zero_8__2__sv2v_reg ;
  assign \xz.mem_with_zero_8__1_  = \xz.mem_with_zero_8__1__sv2v_reg ;
  assign \xz.mem_with_zero_8__0_  = \xz.mem_with_zero_8__0__sv2v_reg ;
  assign \xz.mem_with_zero_7__31_  = \xz.mem_with_zero_7__31__sv2v_reg ;
  assign \xz.mem_with_zero_7__30_  = \xz.mem_with_zero_7__30__sv2v_reg ;
  assign \xz.mem_with_zero_7__29_  = \xz.mem_with_zero_7__29__sv2v_reg ;
  assign \xz.mem_with_zero_7__28_  = \xz.mem_with_zero_7__28__sv2v_reg ;
  assign \xz.mem_with_zero_7__27_  = \xz.mem_with_zero_7__27__sv2v_reg ;
  assign \xz.mem_with_zero_7__26_  = \xz.mem_with_zero_7__26__sv2v_reg ;
  assign \xz.mem_with_zero_7__25_  = \xz.mem_with_zero_7__25__sv2v_reg ;
  assign \xz.mem_with_zero_7__24_  = \xz.mem_with_zero_7__24__sv2v_reg ;
  assign \xz.mem_with_zero_7__23_  = \xz.mem_with_zero_7__23__sv2v_reg ;
  assign \xz.mem_with_zero_7__22_  = \xz.mem_with_zero_7__22__sv2v_reg ;
  assign \xz.mem_with_zero_7__21_  = \xz.mem_with_zero_7__21__sv2v_reg ;
  assign \xz.mem_with_zero_7__20_  = \xz.mem_with_zero_7__20__sv2v_reg ;
  assign \xz.mem_with_zero_7__19_  = \xz.mem_with_zero_7__19__sv2v_reg ;
  assign \xz.mem_with_zero_7__18_  = \xz.mem_with_zero_7__18__sv2v_reg ;
  assign \xz.mem_with_zero_7__17_  = \xz.mem_with_zero_7__17__sv2v_reg ;
  assign \xz.mem_with_zero_7__16_  = \xz.mem_with_zero_7__16__sv2v_reg ;
  assign \xz.mem_with_zero_7__15_  = \xz.mem_with_zero_7__15__sv2v_reg ;
  assign \xz.mem_with_zero_7__14_  = \xz.mem_with_zero_7__14__sv2v_reg ;
  assign \xz.mem_with_zero_7__13_  = \xz.mem_with_zero_7__13__sv2v_reg ;
  assign \xz.mem_with_zero_7__12_  = \xz.mem_with_zero_7__12__sv2v_reg ;
  assign \xz.mem_with_zero_7__11_  = \xz.mem_with_zero_7__11__sv2v_reg ;
  assign \xz.mem_with_zero_7__10_  = \xz.mem_with_zero_7__10__sv2v_reg ;
  assign \xz.mem_with_zero_7__9_  = \xz.mem_with_zero_7__9__sv2v_reg ;
  assign \xz.mem_with_zero_7__8_  = \xz.mem_with_zero_7__8__sv2v_reg ;
  assign \xz.mem_with_zero_7__7_  = \xz.mem_with_zero_7__7__sv2v_reg ;
  assign \xz.mem_with_zero_7__6_  = \xz.mem_with_zero_7__6__sv2v_reg ;
  assign \xz.mem_with_zero_7__5_  = \xz.mem_with_zero_7__5__sv2v_reg ;
  assign \xz.mem_with_zero_7__4_  = \xz.mem_with_zero_7__4__sv2v_reg ;
  assign \xz.mem_with_zero_7__3_  = \xz.mem_with_zero_7__3__sv2v_reg ;
  assign \xz.mem_with_zero_7__2_  = \xz.mem_with_zero_7__2__sv2v_reg ;
  assign \xz.mem_with_zero_7__1_  = \xz.mem_with_zero_7__1__sv2v_reg ;
  assign \xz.mem_with_zero_7__0_  = \xz.mem_with_zero_7__0__sv2v_reg ;
  assign \xz.mem_with_zero_6__31_  = \xz.mem_with_zero_6__31__sv2v_reg ;
  assign \xz.mem_with_zero_6__30_  = \xz.mem_with_zero_6__30__sv2v_reg ;
  assign \xz.mem_with_zero_6__29_  = \xz.mem_with_zero_6__29__sv2v_reg ;
  assign \xz.mem_with_zero_6__28_  = \xz.mem_with_zero_6__28__sv2v_reg ;
  assign \xz.mem_with_zero_6__27_  = \xz.mem_with_zero_6__27__sv2v_reg ;
  assign \xz.mem_with_zero_6__26_  = \xz.mem_with_zero_6__26__sv2v_reg ;
  assign \xz.mem_with_zero_6__25_  = \xz.mem_with_zero_6__25__sv2v_reg ;
  assign \xz.mem_with_zero_6__24_  = \xz.mem_with_zero_6__24__sv2v_reg ;
  assign \xz.mem_with_zero_6__23_  = \xz.mem_with_zero_6__23__sv2v_reg ;
  assign \xz.mem_with_zero_6__22_  = \xz.mem_with_zero_6__22__sv2v_reg ;
  assign \xz.mem_with_zero_6__21_  = \xz.mem_with_zero_6__21__sv2v_reg ;
  assign \xz.mem_with_zero_6__20_  = \xz.mem_with_zero_6__20__sv2v_reg ;
  assign \xz.mem_with_zero_6__19_  = \xz.mem_with_zero_6__19__sv2v_reg ;
  assign \xz.mem_with_zero_6__18_  = \xz.mem_with_zero_6__18__sv2v_reg ;
  assign \xz.mem_with_zero_6__17_  = \xz.mem_with_zero_6__17__sv2v_reg ;
  assign \xz.mem_with_zero_6__16_  = \xz.mem_with_zero_6__16__sv2v_reg ;
  assign \xz.mem_with_zero_6__15_  = \xz.mem_with_zero_6__15__sv2v_reg ;
  assign \xz.mem_with_zero_6__14_  = \xz.mem_with_zero_6__14__sv2v_reg ;
  assign \xz.mem_with_zero_6__13_  = \xz.mem_with_zero_6__13__sv2v_reg ;
  assign \xz.mem_with_zero_6__12_  = \xz.mem_with_zero_6__12__sv2v_reg ;
  assign \xz.mem_with_zero_6__11_  = \xz.mem_with_zero_6__11__sv2v_reg ;
  assign \xz.mem_with_zero_6__10_  = \xz.mem_with_zero_6__10__sv2v_reg ;
  assign \xz.mem_with_zero_6__9_  = \xz.mem_with_zero_6__9__sv2v_reg ;
  assign \xz.mem_with_zero_6__8_  = \xz.mem_with_zero_6__8__sv2v_reg ;
  assign \xz.mem_with_zero_6__7_  = \xz.mem_with_zero_6__7__sv2v_reg ;
  assign \xz.mem_with_zero_6__6_  = \xz.mem_with_zero_6__6__sv2v_reg ;
  assign \xz.mem_with_zero_6__5_  = \xz.mem_with_zero_6__5__sv2v_reg ;
  assign \xz.mem_with_zero_6__4_  = \xz.mem_with_zero_6__4__sv2v_reg ;
  assign \xz.mem_with_zero_6__3_  = \xz.mem_with_zero_6__3__sv2v_reg ;
  assign \xz.mem_with_zero_6__2_  = \xz.mem_with_zero_6__2__sv2v_reg ;
  assign \xz.mem_with_zero_6__1_  = \xz.mem_with_zero_6__1__sv2v_reg ;
  assign \xz.mem_with_zero_6__0_  = \xz.mem_with_zero_6__0__sv2v_reg ;
  assign \xz.mem_with_zero_5__31_  = \xz.mem_with_zero_5__31__sv2v_reg ;
  assign \xz.mem_with_zero_5__30_  = \xz.mem_with_zero_5__30__sv2v_reg ;
  assign \xz.mem_with_zero_5__29_  = \xz.mem_with_zero_5__29__sv2v_reg ;
  assign \xz.mem_with_zero_5__28_  = \xz.mem_with_zero_5__28__sv2v_reg ;
  assign \xz.mem_with_zero_5__27_  = \xz.mem_with_zero_5__27__sv2v_reg ;
  assign \xz.mem_with_zero_5__26_  = \xz.mem_with_zero_5__26__sv2v_reg ;
  assign \xz.mem_with_zero_5__25_  = \xz.mem_with_zero_5__25__sv2v_reg ;
  assign \xz.mem_with_zero_5__24_  = \xz.mem_with_zero_5__24__sv2v_reg ;
  assign \xz.mem_with_zero_5__23_  = \xz.mem_with_zero_5__23__sv2v_reg ;
  assign \xz.mem_with_zero_5__22_  = \xz.mem_with_zero_5__22__sv2v_reg ;
  assign \xz.mem_with_zero_5__21_  = \xz.mem_with_zero_5__21__sv2v_reg ;
  assign \xz.mem_with_zero_5__20_  = \xz.mem_with_zero_5__20__sv2v_reg ;
  assign \xz.mem_with_zero_5__19_  = \xz.mem_with_zero_5__19__sv2v_reg ;
  assign \xz.mem_with_zero_5__18_  = \xz.mem_with_zero_5__18__sv2v_reg ;
  assign \xz.mem_with_zero_5__17_  = \xz.mem_with_zero_5__17__sv2v_reg ;
  assign \xz.mem_with_zero_5__16_  = \xz.mem_with_zero_5__16__sv2v_reg ;
  assign \xz.mem_with_zero_5__15_  = \xz.mem_with_zero_5__15__sv2v_reg ;
  assign \xz.mem_with_zero_5__14_  = \xz.mem_with_zero_5__14__sv2v_reg ;
  assign \xz.mem_with_zero_5__13_  = \xz.mem_with_zero_5__13__sv2v_reg ;
  assign \xz.mem_with_zero_5__12_  = \xz.mem_with_zero_5__12__sv2v_reg ;
  assign \xz.mem_with_zero_5__11_  = \xz.mem_with_zero_5__11__sv2v_reg ;
  assign \xz.mem_with_zero_5__10_  = \xz.mem_with_zero_5__10__sv2v_reg ;
  assign \xz.mem_with_zero_5__9_  = \xz.mem_with_zero_5__9__sv2v_reg ;
  assign \xz.mem_with_zero_5__8_  = \xz.mem_with_zero_5__8__sv2v_reg ;
  assign \xz.mem_with_zero_5__7_  = \xz.mem_with_zero_5__7__sv2v_reg ;
  assign \xz.mem_with_zero_5__6_  = \xz.mem_with_zero_5__6__sv2v_reg ;
  assign \xz.mem_with_zero_5__5_  = \xz.mem_with_zero_5__5__sv2v_reg ;
  assign \xz.mem_with_zero_5__4_  = \xz.mem_with_zero_5__4__sv2v_reg ;
  assign \xz.mem_with_zero_5__3_  = \xz.mem_with_zero_5__3__sv2v_reg ;
  assign \xz.mem_with_zero_5__2_  = \xz.mem_with_zero_5__2__sv2v_reg ;
  assign \xz.mem_with_zero_5__1_  = \xz.mem_with_zero_5__1__sv2v_reg ;
  assign \xz.mem_with_zero_5__0_  = \xz.mem_with_zero_5__0__sv2v_reg ;
  assign \xz.mem_with_zero_4__31_  = \xz.mem_with_zero_4__31__sv2v_reg ;
  assign \xz.mem_with_zero_4__30_  = \xz.mem_with_zero_4__30__sv2v_reg ;
  assign \xz.mem_with_zero_4__29_  = \xz.mem_with_zero_4__29__sv2v_reg ;
  assign \xz.mem_with_zero_4__28_  = \xz.mem_with_zero_4__28__sv2v_reg ;
  assign \xz.mem_with_zero_4__27_  = \xz.mem_with_zero_4__27__sv2v_reg ;
  assign \xz.mem_with_zero_4__26_  = \xz.mem_with_zero_4__26__sv2v_reg ;
  assign \xz.mem_with_zero_4__25_  = \xz.mem_with_zero_4__25__sv2v_reg ;
  assign \xz.mem_with_zero_4__24_  = \xz.mem_with_zero_4__24__sv2v_reg ;
  assign \xz.mem_with_zero_4__23_  = \xz.mem_with_zero_4__23__sv2v_reg ;
  assign \xz.mem_with_zero_4__22_  = \xz.mem_with_zero_4__22__sv2v_reg ;
  assign \xz.mem_with_zero_4__21_  = \xz.mem_with_zero_4__21__sv2v_reg ;
  assign \xz.mem_with_zero_4__20_  = \xz.mem_with_zero_4__20__sv2v_reg ;
  assign \xz.mem_with_zero_4__19_  = \xz.mem_with_zero_4__19__sv2v_reg ;
  assign \xz.mem_with_zero_4__18_  = \xz.mem_with_zero_4__18__sv2v_reg ;
  assign \xz.mem_with_zero_4__17_  = \xz.mem_with_zero_4__17__sv2v_reg ;
  assign \xz.mem_with_zero_4__16_  = \xz.mem_with_zero_4__16__sv2v_reg ;
  assign \xz.mem_with_zero_4__15_  = \xz.mem_with_zero_4__15__sv2v_reg ;
  assign \xz.mem_with_zero_4__14_  = \xz.mem_with_zero_4__14__sv2v_reg ;
  assign \xz.mem_with_zero_4__13_  = \xz.mem_with_zero_4__13__sv2v_reg ;
  assign \xz.mem_with_zero_4__12_  = \xz.mem_with_zero_4__12__sv2v_reg ;
  assign \xz.mem_with_zero_4__11_  = \xz.mem_with_zero_4__11__sv2v_reg ;
  assign \xz.mem_with_zero_4__10_  = \xz.mem_with_zero_4__10__sv2v_reg ;
  assign \xz.mem_with_zero_4__9_  = \xz.mem_with_zero_4__9__sv2v_reg ;
  assign \xz.mem_with_zero_4__8_  = \xz.mem_with_zero_4__8__sv2v_reg ;
  assign \xz.mem_with_zero_4__7_  = \xz.mem_with_zero_4__7__sv2v_reg ;
  assign \xz.mem_with_zero_4__6_  = \xz.mem_with_zero_4__6__sv2v_reg ;
  assign \xz.mem_with_zero_4__5_  = \xz.mem_with_zero_4__5__sv2v_reg ;
  assign \xz.mem_with_zero_4__4_  = \xz.mem_with_zero_4__4__sv2v_reg ;
  assign \xz.mem_with_zero_4__3_  = \xz.mem_with_zero_4__3__sv2v_reg ;
  assign \xz.mem_with_zero_4__2_  = \xz.mem_with_zero_4__2__sv2v_reg ;
  assign \xz.mem_with_zero_4__1_  = \xz.mem_with_zero_4__1__sv2v_reg ;
  assign \xz.mem_with_zero_4__0_  = \xz.mem_with_zero_4__0__sv2v_reg ;
  assign \xz.mem_with_zero_3__31_  = \xz.mem_with_zero_3__31__sv2v_reg ;
  assign \xz.mem_with_zero_3__30_  = \xz.mem_with_zero_3__30__sv2v_reg ;
  assign \xz.mem_with_zero_3__29_  = \xz.mem_with_zero_3__29__sv2v_reg ;
  assign \xz.mem_with_zero_3__28_  = \xz.mem_with_zero_3__28__sv2v_reg ;
  assign \xz.mem_with_zero_3__27_  = \xz.mem_with_zero_3__27__sv2v_reg ;
  assign \xz.mem_with_zero_3__26_  = \xz.mem_with_zero_3__26__sv2v_reg ;
  assign \xz.mem_with_zero_3__25_  = \xz.mem_with_zero_3__25__sv2v_reg ;
  assign \xz.mem_with_zero_3__24_  = \xz.mem_with_zero_3__24__sv2v_reg ;
  assign \xz.mem_with_zero_3__23_  = \xz.mem_with_zero_3__23__sv2v_reg ;
  assign \xz.mem_with_zero_3__22_  = \xz.mem_with_zero_3__22__sv2v_reg ;
  assign \xz.mem_with_zero_3__21_  = \xz.mem_with_zero_3__21__sv2v_reg ;
  assign \xz.mem_with_zero_3__20_  = \xz.mem_with_zero_3__20__sv2v_reg ;
  assign \xz.mem_with_zero_3__19_  = \xz.mem_with_zero_3__19__sv2v_reg ;
  assign \xz.mem_with_zero_3__18_  = \xz.mem_with_zero_3__18__sv2v_reg ;
  assign \xz.mem_with_zero_3__17_  = \xz.mem_with_zero_3__17__sv2v_reg ;
  assign \xz.mem_with_zero_3__16_  = \xz.mem_with_zero_3__16__sv2v_reg ;
  assign \xz.mem_with_zero_3__15_  = \xz.mem_with_zero_3__15__sv2v_reg ;
  assign \xz.mem_with_zero_3__14_  = \xz.mem_with_zero_3__14__sv2v_reg ;
  assign \xz.mem_with_zero_3__13_  = \xz.mem_with_zero_3__13__sv2v_reg ;
  assign \xz.mem_with_zero_3__12_  = \xz.mem_with_zero_3__12__sv2v_reg ;
  assign \xz.mem_with_zero_3__11_  = \xz.mem_with_zero_3__11__sv2v_reg ;
  assign \xz.mem_with_zero_3__10_  = \xz.mem_with_zero_3__10__sv2v_reg ;
  assign \xz.mem_with_zero_3__9_  = \xz.mem_with_zero_3__9__sv2v_reg ;
  assign \xz.mem_with_zero_3__8_  = \xz.mem_with_zero_3__8__sv2v_reg ;
  assign \xz.mem_with_zero_3__7_  = \xz.mem_with_zero_3__7__sv2v_reg ;
  assign \xz.mem_with_zero_3__6_  = \xz.mem_with_zero_3__6__sv2v_reg ;
  assign \xz.mem_with_zero_3__5_  = \xz.mem_with_zero_3__5__sv2v_reg ;
  assign \xz.mem_with_zero_3__4_  = \xz.mem_with_zero_3__4__sv2v_reg ;
  assign \xz.mem_with_zero_3__3_  = \xz.mem_with_zero_3__3__sv2v_reg ;
  assign \xz.mem_with_zero_3__2_  = \xz.mem_with_zero_3__2__sv2v_reg ;
  assign \xz.mem_with_zero_3__1_  = \xz.mem_with_zero_3__1__sv2v_reg ;
  assign \xz.mem_with_zero_3__0_  = \xz.mem_with_zero_3__0__sv2v_reg ;
  assign \xz.mem_with_zero_2__31_  = \xz.mem_with_zero_2__31__sv2v_reg ;
  assign \xz.mem_with_zero_2__30_  = \xz.mem_with_zero_2__30__sv2v_reg ;
  assign \xz.mem_with_zero_2__29_  = \xz.mem_with_zero_2__29__sv2v_reg ;
  assign \xz.mem_with_zero_2__28_  = \xz.mem_with_zero_2__28__sv2v_reg ;
  assign \xz.mem_with_zero_2__27_  = \xz.mem_with_zero_2__27__sv2v_reg ;
  assign \xz.mem_with_zero_2__26_  = \xz.mem_with_zero_2__26__sv2v_reg ;
  assign \xz.mem_with_zero_2__25_  = \xz.mem_with_zero_2__25__sv2v_reg ;
  assign \xz.mem_with_zero_2__24_  = \xz.mem_with_zero_2__24__sv2v_reg ;
  assign \xz.mem_with_zero_2__23_  = \xz.mem_with_zero_2__23__sv2v_reg ;
  assign \xz.mem_with_zero_2__22_  = \xz.mem_with_zero_2__22__sv2v_reg ;
  assign \xz.mem_with_zero_2__21_  = \xz.mem_with_zero_2__21__sv2v_reg ;
  assign \xz.mem_with_zero_2__20_  = \xz.mem_with_zero_2__20__sv2v_reg ;
  assign \xz.mem_with_zero_2__19_  = \xz.mem_with_zero_2__19__sv2v_reg ;
  assign \xz.mem_with_zero_2__18_  = \xz.mem_with_zero_2__18__sv2v_reg ;
  assign \xz.mem_with_zero_2__17_  = \xz.mem_with_zero_2__17__sv2v_reg ;
  assign \xz.mem_with_zero_2__16_  = \xz.mem_with_zero_2__16__sv2v_reg ;
  assign \xz.mem_with_zero_2__15_  = \xz.mem_with_zero_2__15__sv2v_reg ;
  assign \xz.mem_with_zero_2__14_  = \xz.mem_with_zero_2__14__sv2v_reg ;
  assign \xz.mem_with_zero_2__13_  = \xz.mem_with_zero_2__13__sv2v_reg ;
  assign \xz.mem_with_zero_2__12_  = \xz.mem_with_zero_2__12__sv2v_reg ;
  assign \xz.mem_with_zero_2__11_  = \xz.mem_with_zero_2__11__sv2v_reg ;
  assign \xz.mem_with_zero_2__10_  = \xz.mem_with_zero_2__10__sv2v_reg ;
  assign \xz.mem_with_zero_2__9_  = \xz.mem_with_zero_2__9__sv2v_reg ;
  assign \xz.mem_with_zero_2__8_  = \xz.mem_with_zero_2__8__sv2v_reg ;
  assign \xz.mem_with_zero_2__7_  = \xz.mem_with_zero_2__7__sv2v_reg ;
  assign \xz.mem_with_zero_2__6_  = \xz.mem_with_zero_2__6__sv2v_reg ;
  assign \xz.mem_with_zero_2__5_  = \xz.mem_with_zero_2__5__sv2v_reg ;
  assign \xz.mem_with_zero_2__4_  = \xz.mem_with_zero_2__4__sv2v_reg ;
  assign \xz.mem_with_zero_2__3_  = \xz.mem_with_zero_2__3__sv2v_reg ;
  assign \xz.mem_with_zero_2__2_  = \xz.mem_with_zero_2__2__sv2v_reg ;
  assign \xz.mem_with_zero_2__1_  = \xz.mem_with_zero_2__1__sv2v_reg ;
  assign \xz.mem_with_zero_2__0_  = \xz.mem_with_zero_2__0__sv2v_reg ;
  assign \xz.mem_with_zero_1__31_  = \xz.mem_with_zero_1__31__sv2v_reg ;
  assign \xz.mem_with_zero_1__30_  = \xz.mem_with_zero_1__30__sv2v_reg ;
  assign \xz.mem_with_zero_1__29_  = \xz.mem_with_zero_1__29__sv2v_reg ;
  assign \xz.mem_with_zero_1__28_  = \xz.mem_with_zero_1__28__sv2v_reg ;
  assign \xz.mem_with_zero_1__27_  = \xz.mem_with_zero_1__27__sv2v_reg ;
  assign \xz.mem_with_zero_1__26_  = \xz.mem_with_zero_1__26__sv2v_reg ;
  assign \xz.mem_with_zero_1__25_  = \xz.mem_with_zero_1__25__sv2v_reg ;
  assign \xz.mem_with_zero_1__24_  = \xz.mem_with_zero_1__24__sv2v_reg ;
  assign \xz.mem_with_zero_1__23_  = \xz.mem_with_zero_1__23__sv2v_reg ;
  assign \xz.mem_with_zero_1__22_  = \xz.mem_with_zero_1__22__sv2v_reg ;
  assign \xz.mem_with_zero_1__21_  = \xz.mem_with_zero_1__21__sv2v_reg ;
  assign \xz.mem_with_zero_1__20_  = \xz.mem_with_zero_1__20__sv2v_reg ;
  assign \xz.mem_with_zero_1__19_  = \xz.mem_with_zero_1__19__sv2v_reg ;
  assign \xz.mem_with_zero_1__18_  = \xz.mem_with_zero_1__18__sv2v_reg ;
  assign \xz.mem_with_zero_1__17_  = \xz.mem_with_zero_1__17__sv2v_reg ;
  assign \xz.mem_with_zero_1__16_  = \xz.mem_with_zero_1__16__sv2v_reg ;
  assign \xz.mem_with_zero_1__15_  = \xz.mem_with_zero_1__15__sv2v_reg ;
  assign \xz.mem_with_zero_1__14_  = \xz.mem_with_zero_1__14__sv2v_reg ;
  assign \xz.mem_with_zero_1__13_  = \xz.mem_with_zero_1__13__sv2v_reg ;
  assign \xz.mem_with_zero_1__12_  = \xz.mem_with_zero_1__12__sv2v_reg ;
  assign \xz.mem_with_zero_1__11_  = \xz.mem_with_zero_1__11__sv2v_reg ;
  assign \xz.mem_with_zero_1__10_  = \xz.mem_with_zero_1__10__sv2v_reg ;
  assign \xz.mem_with_zero_1__9_  = \xz.mem_with_zero_1__9__sv2v_reg ;
  assign \xz.mem_with_zero_1__8_  = \xz.mem_with_zero_1__8__sv2v_reg ;
  assign \xz.mem_with_zero_1__7_  = \xz.mem_with_zero_1__7__sv2v_reg ;
  assign \xz.mem_with_zero_1__6_  = \xz.mem_with_zero_1__6__sv2v_reg ;
  assign \xz.mem_with_zero_1__5_  = \xz.mem_with_zero_1__5__sv2v_reg ;
  assign \xz.mem_with_zero_1__4_  = \xz.mem_with_zero_1__4__sv2v_reg ;
  assign \xz.mem_with_zero_1__3_  = \xz.mem_with_zero_1__3__sv2v_reg ;
  assign \xz.mem_with_zero_1__2_  = \xz.mem_with_zero_1__2__sv2v_reg ;
  assign \xz.mem_with_zero_1__1_  = \xz.mem_with_zero_1__1__sv2v_reg ;
  assign \xz.mem_with_zero_1__0_  = \xz.mem_with_zero_1__0__sv2v_reg ;
  assign r_data_o[31] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__31_  : 
                        (N46)? \xz.mem_with_zero_2__31_  : 
                        (N48)? \xz.mem_with_zero_3__31_  : 
                        (N50)? \xz.mem_with_zero_4__31_  : 
                        (N52)? \xz.mem_with_zero_5__31_  : 
                        (N54)? \xz.mem_with_zero_6__31_  : 
                        (N56)? \xz.mem_with_zero_7__31_  : 
                        (N58)? \xz.mem_with_zero_8__31_  : 
                        (N60)? \xz.mem_with_zero_9__31_  : 
                        (N62)? \xz.mem_with_zero_10__31_  : 
                        (N64)? \xz.mem_with_zero_11__31_  : 
                        (N66)? \xz.mem_with_zero_12__31_  : 
                        (N68)? \xz.mem_with_zero_13__31_  : 
                        (N70)? \xz.mem_with_zero_14__31_  : 
                        (N72)? \xz.mem_with_zero_15__31_  : 
                        (N43)? \xz.mem_with_zero_16__31_  : 
                        (N45)? \xz.mem_with_zero_17__31_  : 
                        (N47)? \xz.mem_with_zero_18__31_  : 
                        (N49)? \xz.mem_with_zero_19__31_  : 
                        (N51)? \xz.mem_with_zero_20__31_  : 
                        (N53)? \xz.mem_with_zero_21__31_  : 
                        (N55)? \xz.mem_with_zero_22__31_  : 
                        (N57)? \xz.mem_with_zero_23__31_  : 
                        (N59)? \xz.mem_with_zero_24__31_  : 
                        (N61)? \xz.mem_with_zero_25__31_  : 
                        (N63)? \xz.mem_with_zero_26__31_  : 
                        (N65)? \xz.mem_with_zero_27__31_  : 
                        (N67)? \xz.mem_with_zero_28__31_  : 
                        (N69)? \xz.mem_with_zero_29__31_  : 
                        (N71)? \xz.mem_with_zero_30__31_  : 
                        (N73)? \xz.mem_with_zero_31__31_  : 1'b0;
  assign r_data_o[30] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__30_  : 
                        (N46)? \xz.mem_with_zero_2__30_  : 
                        (N48)? \xz.mem_with_zero_3__30_  : 
                        (N50)? \xz.mem_with_zero_4__30_  : 
                        (N52)? \xz.mem_with_zero_5__30_  : 
                        (N54)? \xz.mem_with_zero_6__30_  : 
                        (N56)? \xz.mem_with_zero_7__30_  : 
                        (N58)? \xz.mem_with_zero_8__30_  : 
                        (N60)? \xz.mem_with_zero_9__30_  : 
                        (N62)? \xz.mem_with_zero_10__30_  : 
                        (N64)? \xz.mem_with_zero_11__30_  : 
                        (N66)? \xz.mem_with_zero_12__30_  : 
                        (N68)? \xz.mem_with_zero_13__30_  : 
                        (N70)? \xz.mem_with_zero_14__30_  : 
                        (N72)? \xz.mem_with_zero_15__30_  : 
                        (N43)? \xz.mem_with_zero_16__30_  : 
                        (N45)? \xz.mem_with_zero_17__30_  : 
                        (N47)? \xz.mem_with_zero_18__30_  : 
                        (N49)? \xz.mem_with_zero_19__30_  : 
                        (N51)? \xz.mem_with_zero_20__30_  : 
                        (N53)? \xz.mem_with_zero_21__30_  : 
                        (N55)? \xz.mem_with_zero_22__30_  : 
                        (N57)? \xz.mem_with_zero_23__30_  : 
                        (N59)? \xz.mem_with_zero_24__30_  : 
                        (N61)? \xz.mem_with_zero_25__30_  : 
                        (N63)? \xz.mem_with_zero_26__30_  : 
                        (N65)? \xz.mem_with_zero_27__30_  : 
                        (N67)? \xz.mem_with_zero_28__30_  : 
                        (N69)? \xz.mem_with_zero_29__30_  : 
                        (N71)? \xz.mem_with_zero_30__30_  : 
                        (N73)? \xz.mem_with_zero_31__30_  : 1'b0;
  assign r_data_o[29] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__29_  : 
                        (N46)? \xz.mem_with_zero_2__29_  : 
                        (N48)? \xz.mem_with_zero_3__29_  : 
                        (N50)? \xz.mem_with_zero_4__29_  : 
                        (N52)? \xz.mem_with_zero_5__29_  : 
                        (N54)? \xz.mem_with_zero_6__29_  : 
                        (N56)? \xz.mem_with_zero_7__29_  : 
                        (N58)? \xz.mem_with_zero_8__29_  : 
                        (N60)? \xz.mem_with_zero_9__29_  : 
                        (N62)? \xz.mem_with_zero_10__29_  : 
                        (N64)? \xz.mem_with_zero_11__29_  : 
                        (N66)? \xz.mem_with_zero_12__29_  : 
                        (N68)? \xz.mem_with_zero_13__29_  : 
                        (N70)? \xz.mem_with_zero_14__29_  : 
                        (N72)? \xz.mem_with_zero_15__29_  : 
                        (N43)? \xz.mem_with_zero_16__29_  : 
                        (N45)? \xz.mem_with_zero_17__29_  : 
                        (N47)? \xz.mem_with_zero_18__29_  : 
                        (N49)? \xz.mem_with_zero_19__29_  : 
                        (N51)? \xz.mem_with_zero_20__29_  : 
                        (N53)? \xz.mem_with_zero_21__29_  : 
                        (N55)? \xz.mem_with_zero_22__29_  : 
                        (N57)? \xz.mem_with_zero_23__29_  : 
                        (N59)? \xz.mem_with_zero_24__29_  : 
                        (N61)? \xz.mem_with_zero_25__29_  : 
                        (N63)? \xz.mem_with_zero_26__29_  : 
                        (N65)? \xz.mem_with_zero_27__29_  : 
                        (N67)? \xz.mem_with_zero_28__29_  : 
                        (N69)? \xz.mem_with_zero_29__29_  : 
                        (N71)? \xz.mem_with_zero_30__29_  : 
                        (N73)? \xz.mem_with_zero_31__29_  : 1'b0;
  assign r_data_o[28] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__28_  : 
                        (N46)? \xz.mem_with_zero_2__28_  : 
                        (N48)? \xz.mem_with_zero_3__28_  : 
                        (N50)? \xz.mem_with_zero_4__28_  : 
                        (N52)? \xz.mem_with_zero_5__28_  : 
                        (N54)? \xz.mem_with_zero_6__28_  : 
                        (N56)? \xz.mem_with_zero_7__28_  : 
                        (N58)? \xz.mem_with_zero_8__28_  : 
                        (N60)? \xz.mem_with_zero_9__28_  : 
                        (N62)? \xz.mem_with_zero_10__28_  : 
                        (N64)? \xz.mem_with_zero_11__28_  : 
                        (N66)? \xz.mem_with_zero_12__28_  : 
                        (N68)? \xz.mem_with_zero_13__28_  : 
                        (N70)? \xz.mem_with_zero_14__28_  : 
                        (N72)? \xz.mem_with_zero_15__28_  : 
                        (N43)? \xz.mem_with_zero_16__28_  : 
                        (N45)? \xz.mem_with_zero_17__28_  : 
                        (N47)? \xz.mem_with_zero_18__28_  : 
                        (N49)? \xz.mem_with_zero_19__28_  : 
                        (N51)? \xz.mem_with_zero_20__28_  : 
                        (N53)? \xz.mem_with_zero_21__28_  : 
                        (N55)? \xz.mem_with_zero_22__28_  : 
                        (N57)? \xz.mem_with_zero_23__28_  : 
                        (N59)? \xz.mem_with_zero_24__28_  : 
                        (N61)? \xz.mem_with_zero_25__28_  : 
                        (N63)? \xz.mem_with_zero_26__28_  : 
                        (N65)? \xz.mem_with_zero_27__28_  : 
                        (N67)? \xz.mem_with_zero_28__28_  : 
                        (N69)? \xz.mem_with_zero_29__28_  : 
                        (N71)? \xz.mem_with_zero_30__28_  : 
                        (N73)? \xz.mem_with_zero_31__28_  : 1'b0;
  assign r_data_o[27] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__27_  : 
                        (N46)? \xz.mem_with_zero_2__27_  : 
                        (N48)? \xz.mem_with_zero_3__27_  : 
                        (N50)? \xz.mem_with_zero_4__27_  : 
                        (N52)? \xz.mem_with_zero_5__27_  : 
                        (N54)? \xz.mem_with_zero_6__27_  : 
                        (N56)? \xz.mem_with_zero_7__27_  : 
                        (N58)? \xz.mem_with_zero_8__27_  : 
                        (N60)? \xz.mem_with_zero_9__27_  : 
                        (N62)? \xz.mem_with_zero_10__27_  : 
                        (N64)? \xz.mem_with_zero_11__27_  : 
                        (N66)? \xz.mem_with_zero_12__27_  : 
                        (N68)? \xz.mem_with_zero_13__27_  : 
                        (N70)? \xz.mem_with_zero_14__27_  : 
                        (N72)? \xz.mem_with_zero_15__27_  : 
                        (N43)? \xz.mem_with_zero_16__27_  : 
                        (N45)? \xz.mem_with_zero_17__27_  : 
                        (N47)? \xz.mem_with_zero_18__27_  : 
                        (N49)? \xz.mem_with_zero_19__27_  : 
                        (N51)? \xz.mem_with_zero_20__27_  : 
                        (N53)? \xz.mem_with_zero_21__27_  : 
                        (N55)? \xz.mem_with_zero_22__27_  : 
                        (N57)? \xz.mem_with_zero_23__27_  : 
                        (N59)? \xz.mem_with_zero_24__27_  : 
                        (N61)? \xz.mem_with_zero_25__27_  : 
                        (N63)? \xz.mem_with_zero_26__27_  : 
                        (N65)? \xz.mem_with_zero_27__27_  : 
                        (N67)? \xz.mem_with_zero_28__27_  : 
                        (N69)? \xz.mem_with_zero_29__27_  : 
                        (N71)? \xz.mem_with_zero_30__27_  : 
                        (N73)? \xz.mem_with_zero_31__27_  : 1'b0;
  assign r_data_o[26] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__26_  : 
                        (N46)? \xz.mem_with_zero_2__26_  : 
                        (N48)? \xz.mem_with_zero_3__26_  : 
                        (N50)? \xz.mem_with_zero_4__26_  : 
                        (N52)? \xz.mem_with_zero_5__26_  : 
                        (N54)? \xz.mem_with_zero_6__26_  : 
                        (N56)? \xz.mem_with_zero_7__26_  : 
                        (N58)? \xz.mem_with_zero_8__26_  : 
                        (N60)? \xz.mem_with_zero_9__26_  : 
                        (N62)? \xz.mem_with_zero_10__26_  : 
                        (N64)? \xz.mem_with_zero_11__26_  : 
                        (N66)? \xz.mem_with_zero_12__26_  : 
                        (N68)? \xz.mem_with_zero_13__26_  : 
                        (N70)? \xz.mem_with_zero_14__26_  : 
                        (N72)? \xz.mem_with_zero_15__26_  : 
                        (N43)? \xz.mem_with_zero_16__26_  : 
                        (N45)? \xz.mem_with_zero_17__26_  : 
                        (N47)? \xz.mem_with_zero_18__26_  : 
                        (N49)? \xz.mem_with_zero_19__26_  : 
                        (N51)? \xz.mem_with_zero_20__26_  : 
                        (N53)? \xz.mem_with_zero_21__26_  : 
                        (N55)? \xz.mem_with_zero_22__26_  : 
                        (N57)? \xz.mem_with_zero_23__26_  : 
                        (N59)? \xz.mem_with_zero_24__26_  : 
                        (N61)? \xz.mem_with_zero_25__26_  : 
                        (N63)? \xz.mem_with_zero_26__26_  : 
                        (N65)? \xz.mem_with_zero_27__26_  : 
                        (N67)? \xz.mem_with_zero_28__26_  : 
                        (N69)? \xz.mem_with_zero_29__26_  : 
                        (N71)? \xz.mem_with_zero_30__26_  : 
                        (N73)? \xz.mem_with_zero_31__26_  : 1'b0;
  assign r_data_o[25] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__25_  : 
                        (N46)? \xz.mem_with_zero_2__25_  : 
                        (N48)? \xz.mem_with_zero_3__25_  : 
                        (N50)? \xz.mem_with_zero_4__25_  : 
                        (N52)? \xz.mem_with_zero_5__25_  : 
                        (N54)? \xz.mem_with_zero_6__25_  : 
                        (N56)? \xz.mem_with_zero_7__25_  : 
                        (N58)? \xz.mem_with_zero_8__25_  : 
                        (N60)? \xz.mem_with_zero_9__25_  : 
                        (N62)? \xz.mem_with_zero_10__25_  : 
                        (N64)? \xz.mem_with_zero_11__25_  : 
                        (N66)? \xz.mem_with_zero_12__25_  : 
                        (N68)? \xz.mem_with_zero_13__25_  : 
                        (N70)? \xz.mem_with_zero_14__25_  : 
                        (N72)? \xz.mem_with_zero_15__25_  : 
                        (N43)? \xz.mem_with_zero_16__25_  : 
                        (N45)? \xz.mem_with_zero_17__25_  : 
                        (N47)? \xz.mem_with_zero_18__25_  : 
                        (N49)? \xz.mem_with_zero_19__25_  : 
                        (N51)? \xz.mem_with_zero_20__25_  : 
                        (N53)? \xz.mem_with_zero_21__25_  : 
                        (N55)? \xz.mem_with_zero_22__25_  : 
                        (N57)? \xz.mem_with_zero_23__25_  : 
                        (N59)? \xz.mem_with_zero_24__25_  : 
                        (N61)? \xz.mem_with_zero_25__25_  : 
                        (N63)? \xz.mem_with_zero_26__25_  : 
                        (N65)? \xz.mem_with_zero_27__25_  : 
                        (N67)? \xz.mem_with_zero_28__25_  : 
                        (N69)? \xz.mem_with_zero_29__25_  : 
                        (N71)? \xz.mem_with_zero_30__25_  : 
                        (N73)? \xz.mem_with_zero_31__25_  : 1'b0;
  assign r_data_o[24] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__24_  : 
                        (N46)? \xz.mem_with_zero_2__24_  : 
                        (N48)? \xz.mem_with_zero_3__24_  : 
                        (N50)? \xz.mem_with_zero_4__24_  : 
                        (N52)? \xz.mem_with_zero_5__24_  : 
                        (N54)? \xz.mem_with_zero_6__24_  : 
                        (N56)? \xz.mem_with_zero_7__24_  : 
                        (N58)? \xz.mem_with_zero_8__24_  : 
                        (N60)? \xz.mem_with_zero_9__24_  : 
                        (N62)? \xz.mem_with_zero_10__24_  : 
                        (N64)? \xz.mem_with_zero_11__24_  : 
                        (N66)? \xz.mem_with_zero_12__24_  : 
                        (N68)? \xz.mem_with_zero_13__24_  : 
                        (N70)? \xz.mem_with_zero_14__24_  : 
                        (N72)? \xz.mem_with_zero_15__24_  : 
                        (N43)? \xz.mem_with_zero_16__24_  : 
                        (N45)? \xz.mem_with_zero_17__24_  : 
                        (N47)? \xz.mem_with_zero_18__24_  : 
                        (N49)? \xz.mem_with_zero_19__24_  : 
                        (N51)? \xz.mem_with_zero_20__24_  : 
                        (N53)? \xz.mem_with_zero_21__24_  : 
                        (N55)? \xz.mem_with_zero_22__24_  : 
                        (N57)? \xz.mem_with_zero_23__24_  : 
                        (N59)? \xz.mem_with_zero_24__24_  : 
                        (N61)? \xz.mem_with_zero_25__24_  : 
                        (N63)? \xz.mem_with_zero_26__24_  : 
                        (N65)? \xz.mem_with_zero_27__24_  : 
                        (N67)? \xz.mem_with_zero_28__24_  : 
                        (N69)? \xz.mem_with_zero_29__24_  : 
                        (N71)? \xz.mem_with_zero_30__24_  : 
                        (N73)? \xz.mem_with_zero_31__24_  : 1'b0;
  assign r_data_o[23] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__23_  : 
                        (N46)? \xz.mem_with_zero_2__23_  : 
                        (N48)? \xz.mem_with_zero_3__23_  : 
                        (N50)? \xz.mem_with_zero_4__23_  : 
                        (N52)? \xz.mem_with_zero_5__23_  : 
                        (N54)? \xz.mem_with_zero_6__23_  : 
                        (N56)? \xz.mem_with_zero_7__23_  : 
                        (N58)? \xz.mem_with_zero_8__23_  : 
                        (N60)? \xz.mem_with_zero_9__23_  : 
                        (N62)? \xz.mem_with_zero_10__23_  : 
                        (N64)? \xz.mem_with_zero_11__23_  : 
                        (N66)? \xz.mem_with_zero_12__23_  : 
                        (N68)? \xz.mem_with_zero_13__23_  : 
                        (N70)? \xz.mem_with_zero_14__23_  : 
                        (N72)? \xz.mem_with_zero_15__23_  : 
                        (N43)? \xz.mem_with_zero_16__23_  : 
                        (N45)? \xz.mem_with_zero_17__23_  : 
                        (N47)? \xz.mem_with_zero_18__23_  : 
                        (N49)? \xz.mem_with_zero_19__23_  : 
                        (N51)? \xz.mem_with_zero_20__23_  : 
                        (N53)? \xz.mem_with_zero_21__23_  : 
                        (N55)? \xz.mem_with_zero_22__23_  : 
                        (N57)? \xz.mem_with_zero_23__23_  : 
                        (N59)? \xz.mem_with_zero_24__23_  : 
                        (N61)? \xz.mem_with_zero_25__23_  : 
                        (N63)? \xz.mem_with_zero_26__23_  : 
                        (N65)? \xz.mem_with_zero_27__23_  : 
                        (N67)? \xz.mem_with_zero_28__23_  : 
                        (N69)? \xz.mem_with_zero_29__23_  : 
                        (N71)? \xz.mem_with_zero_30__23_  : 
                        (N73)? \xz.mem_with_zero_31__23_  : 1'b0;
  assign r_data_o[22] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__22_  : 
                        (N46)? \xz.mem_with_zero_2__22_  : 
                        (N48)? \xz.mem_with_zero_3__22_  : 
                        (N50)? \xz.mem_with_zero_4__22_  : 
                        (N52)? \xz.mem_with_zero_5__22_  : 
                        (N54)? \xz.mem_with_zero_6__22_  : 
                        (N56)? \xz.mem_with_zero_7__22_  : 
                        (N58)? \xz.mem_with_zero_8__22_  : 
                        (N60)? \xz.mem_with_zero_9__22_  : 
                        (N62)? \xz.mem_with_zero_10__22_  : 
                        (N64)? \xz.mem_with_zero_11__22_  : 
                        (N66)? \xz.mem_with_zero_12__22_  : 
                        (N68)? \xz.mem_with_zero_13__22_  : 
                        (N70)? \xz.mem_with_zero_14__22_  : 
                        (N72)? \xz.mem_with_zero_15__22_  : 
                        (N43)? \xz.mem_with_zero_16__22_  : 
                        (N45)? \xz.mem_with_zero_17__22_  : 
                        (N47)? \xz.mem_with_zero_18__22_  : 
                        (N49)? \xz.mem_with_zero_19__22_  : 
                        (N51)? \xz.mem_with_zero_20__22_  : 
                        (N53)? \xz.mem_with_zero_21__22_  : 
                        (N55)? \xz.mem_with_zero_22__22_  : 
                        (N57)? \xz.mem_with_zero_23__22_  : 
                        (N59)? \xz.mem_with_zero_24__22_  : 
                        (N61)? \xz.mem_with_zero_25__22_  : 
                        (N63)? \xz.mem_with_zero_26__22_  : 
                        (N65)? \xz.mem_with_zero_27__22_  : 
                        (N67)? \xz.mem_with_zero_28__22_  : 
                        (N69)? \xz.mem_with_zero_29__22_  : 
                        (N71)? \xz.mem_with_zero_30__22_  : 
                        (N73)? \xz.mem_with_zero_31__22_  : 1'b0;
  assign r_data_o[21] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__21_  : 
                        (N46)? \xz.mem_with_zero_2__21_  : 
                        (N48)? \xz.mem_with_zero_3__21_  : 
                        (N50)? \xz.mem_with_zero_4__21_  : 
                        (N52)? \xz.mem_with_zero_5__21_  : 
                        (N54)? \xz.mem_with_zero_6__21_  : 
                        (N56)? \xz.mem_with_zero_7__21_  : 
                        (N58)? \xz.mem_with_zero_8__21_  : 
                        (N60)? \xz.mem_with_zero_9__21_  : 
                        (N62)? \xz.mem_with_zero_10__21_  : 
                        (N64)? \xz.mem_with_zero_11__21_  : 
                        (N66)? \xz.mem_with_zero_12__21_  : 
                        (N68)? \xz.mem_with_zero_13__21_  : 
                        (N70)? \xz.mem_with_zero_14__21_  : 
                        (N72)? \xz.mem_with_zero_15__21_  : 
                        (N43)? \xz.mem_with_zero_16__21_  : 
                        (N45)? \xz.mem_with_zero_17__21_  : 
                        (N47)? \xz.mem_with_zero_18__21_  : 
                        (N49)? \xz.mem_with_zero_19__21_  : 
                        (N51)? \xz.mem_with_zero_20__21_  : 
                        (N53)? \xz.mem_with_zero_21__21_  : 
                        (N55)? \xz.mem_with_zero_22__21_  : 
                        (N57)? \xz.mem_with_zero_23__21_  : 
                        (N59)? \xz.mem_with_zero_24__21_  : 
                        (N61)? \xz.mem_with_zero_25__21_  : 
                        (N63)? \xz.mem_with_zero_26__21_  : 
                        (N65)? \xz.mem_with_zero_27__21_  : 
                        (N67)? \xz.mem_with_zero_28__21_  : 
                        (N69)? \xz.mem_with_zero_29__21_  : 
                        (N71)? \xz.mem_with_zero_30__21_  : 
                        (N73)? \xz.mem_with_zero_31__21_  : 1'b0;
  assign r_data_o[20] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__20_  : 
                        (N46)? \xz.mem_with_zero_2__20_  : 
                        (N48)? \xz.mem_with_zero_3__20_  : 
                        (N50)? \xz.mem_with_zero_4__20_  : 
                        (N52)? \xz.mem_with_zero_5__20_  : 
                        (N54)? \xz.mem_with_zero_6__20_  : 
                        (N56)? \xz.mem_with_zero_7__20_  : 
                        (N58)? \xz.mem_with_zero_8__20_  : 
                        (N60)? \xz.mem_with_zero_9__20_  : 
                        (N62)? \xz.mem_with_zero_10__20_  : 
                        (N64)? \xz.mem_with_zero_11__20_  : 
                        (N66)? \xz.mem_with_zero_12__20_  : 
                        (N68)? \xz.mem_with_zero_13__20_  : 
                        (N70)? \xz.mem_with_zero_14__20_  : 
                        (N72)? \xz.mem_with_zero_15__20_  : 
                        (N43)? \xz.mem_with_zero_16__20_  : 
                        (N45)? \xz.mem_with_zero_17__20_  : 
                        (N47)? \xz.mem_with_zero_18__20_  : 
                        (N49)? \xz.mem_with_zero_19__20_  : 
                        (N51)? \xz.mem_with_zero_20__20_  : 
                        (N53)? \xz.mem_with_zero_21__20_  : 
                        (N55)? \xz.mem_with_zero_22__20_  : 
                        (N57)? \xz.mem_with_zero_23__20_  : 
                        (N59)? \xz.mem_with_zero_24__20_  : 
                        (N61)? \xz.mem_with_zero_25__20_  : 
                        (N63)? \xz.mem_with_zero_26__20_  : 
                        (N65)? \xz.mem_with_zero_27__20_  : 
                        (N67)? \xz.mem_with_zero_28__20_  : 
                        (N69)? \xz.mem_with_zero_29__20_  : 
                        (N71)? \xz.mem_with_zero_30__20_  : 
                        (N73)? \xz.mem_with_zero_31__20_  : 1'b0;
  assign r_data_o[19] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__19_  : 
                        (N46)? \xz.mem_with_zero_2__19_  : 
                        (N48)? \xz.mem_with_zero_3__19_  : 
                        (N50)? \xz.mem_with_zero_4__19_  : 
                        (N52)? \xz.mem_with_zero_5__19_  : 
                        (N54)? \xz.mem_with_zero_6__19_  : 
                        (N56)? \xz.mem_with_zero_7__19_  : 
                        (N58)? \xz.mem_with_zero_8__19_  : 
                        (N60)? \xz.mem_with_zero_9__19_  : 
                        (N62)? \xz.mem_with_zero_10__19_  : 
                        (N64)? \xz.mem_with_zero_11__19_  : 
                        (N66)? \xz.mem_with_zero_12__19_  : 
                        (N68)? \xz.mem_with_zero_13__19_  : 
                        (N70)? \xz.mem_with_zero_14__19_  : 
                        (N72)? \xz.mem_with_zero_15__19_  : 
                        (N43)? \xz.mem_with_zero_16__19_  : 
                        (N45)? \xz.mem_with_zero_17__19_  : 
                        (N47)? \xz.mem_with_zero_18__19_  : 
                        (N49)? \xz.mem_with_zero_19__19_  : 
                        (N51)? \xz.mem_with_zero_20__19_  : 
                        (N53)? \xz.mem_with_zero_21__19_  : 
                        (N55)? \xz.mem_with_zero_22__19_  : 
                        (N57)? \xz.mem_with_zero_23__19_  : 
                        (N59)? \xz.mem_with_zero_24__19_  : 
                        (N61)? \xz.mem_with_zero_25__19_  : 
                        (N63)? \xz.mem_with_zero_26__19_  : 
                        (N65)? \xz.mem_with_zero_27__19_  : 
                        (N67)? \xz.mem_with_zero_28__19_  : 
                        (N69)? \xz.mem_with_zero_29__19_  : 
                        (N71)? \xz.mem_with_zero_30__19_  : 
                        (N73)? \xz.mem_with_zero_31__19_  : 1'b0;
  assign r_data_o[18] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__18_  : 
                        (N46)? \xz.mem_with_zero_2__18_  : 
                        (N48)? \xz.mem_with_zero_3__18_  : 
                        (N50)? \xz.mem_with_zero_4__18_  : 
                        (N52)? \xz.mem_with_zero_5__18_  : 
                        (N54)? \xz.mem_with_zero_6__18_  : 
                        (N56)? \xz.mem_with_zero_7__18_  : 
                        (N58)? \xz.mem_with_zero_8__18_  : 
                        (N60)? \xz.mem_with_zero_9__18_  : 
                        (N62)? \xz.mem_with_zero_10__18_  : 
                        (N64)? \xz.mem_with_zero_11__18_  : 
                        (N66)? \xz.mem_with_zero_12__18_  : 
                        (N68)? \xz.mem_with_zero_13__18_  : 
                        (N70)? \xz.mem_with_zero_14__18_  : 
                        (N72)? \xz.mem_with_zero_15__18_  : 
                        (N43)? \xz.mem_with_zero_16__18_  : 
                        (N45)? \xz.mem_with_zero_17__18_  : 
                        (N47)? \xz.mem_with_zero_18__18_  : 
                        (N49)? \xz.mem_with_zero_19__18_  : 
                        (N51)? \xz.mem_with_zero_20__18_  : 
                        (N53)? \xz.mem_with_zero_21__18_  : 
                        (N55)? \xz.mem_with_zero_22__18_  : 
                        (N57)? \xz.mem_with_zero_23__18_  : 
                        (N59)? \xz.mem_with_zero_24__18_  : 
                        (N61)? \xz.mem_with_zero_25__18_  : 
                        (N63)? \xz.mem_with_zero_26__18_  : 
                        (N65)? \xz.mem_with_zero_27__18_  : 
                        (N67)? \xz.mem_with_zero_28__18_  : 
                        (N69)? \xz.mem_with_zero_29__18_  : 
                        (N71)? \xz.mem_with_zero_30__18_  : 
                        (N73)? \xz.mem_with_zero_31__18_  : 1'b0;
  assign r_data_o[17] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__17_  : 
                        (N46)? \xz.mem_with_zero_2__17_  : 
                        (N48)? \xz.mem_with_zero_3__17_  : 
                        (N50)? \xz.mem_with_zero_4__17_  : 
                        (N52)? \xz.mem_with_zero_5__17_  : 
                        (N54)? \xz.mem_with_zero_6__17_  : 
                        (N56)? \xz.mem_with_zero_7__17_  : 
                        (N58)? \xz.mem_with_zero_8__17_  : 
                        (N60)? \xz.mem_with_zero_9__17_  : 
                        (N62)? \xz.mem_with_zero_10__17_  : 
                        (N64)? \xz.mem_with_zero_11__17_  : 
                        (N66)? \xz.mem_with_zero_12__17_  : 
                        (N68)? \xz.mem_with_zero_13__17_  : 
                        (N70)? \xz.mem_with_zero_14__17_  : 
                        (N72)? \xz.mem_with_zero_15__17_  : 
                        (N43)? \xz.mem_with_zero_16__17_  : 
                        (N45)? \xz.mem_with_zero_17__17_  : 
                        (N47)? \xz.mem_with_zero_18__17_  : 
                        (N49)? \xz.mem_with_zero_19__17_  : 
                        (N51)? \xz.mem_with_zero_20__17_  : 
                        (N53)? \xz.mem_with_zero_21__17_  : 
                        (N55)? \xz.mem_with_zero_22__17_  : 
                        (N57)? \xz.mem_with_zero_23__17_  : 
                        (N59)? \xz.mem_with_zero_24__17_  : 
                        (N61)? \xz.mem_with_zero_25__17_  : 
                        (N63)? \xz.mem_with_zero_26__17_  : 
                        (N65)? \xz.mem_with_zero_27__17_  : 
                        (N67)? \xz.mem_with_zero_28__17_  : 
                        (N69)? \xz.mem_with_zero_29__17_  : 
                        (N71)? \xz.mem_with_zero_30__17_  : 
                        (N73)? \xz.mem_with_zero_31__17_  : 1'b0;
  assign r_data_o[16] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__16_  : 
                        (N46)? \xz.mem_with_zero_2__16_  : 
                        (N48)? \xz.mem_with_zero_3__16_  : 
                        (N50)? \xz.mem_with_zero_4__16_  : 
                        (N52)? \xz.mem_with_zero_5__16_  : 
                        (N54)? \xz.mem_with_zero_6__16_  : 
                        (N56)? \xz.mem_with_zero_7__16_  : 
                        (N58)? \xz.mem_with_zero_8__16_  : 
                        (N60)? \xz.mem_with_zero_9__16_  : 
                        (N62)? \xz.mem_with_zero_10__16_  : 
                        (N64)? \xz.mem_with_zero_11__16_  : 
                        (N66)? \xz.mem_with_zero_12__16_  : 
                        (N68)? \xz.mem_with_zero_13__16_  : 
                        (N70)? \xz.mem_with_zero_14__16_  : 
                        (N72)? \xz.mem_with_zero_15__16_  : 
                        (N43)? \xz.mem_with_zero_16__16_  : 
                        (N45)? \xz.mem_with_zero_17__16_  : 
                        (N47)? \xz.mem_with_zero_18__16_  : 
                        (N49)? \xz.mem_with_zero_19__16_  : 
                        (N51)? \xz.mem_with_zero_20__16_  : 
                        (N53)? \xz.mem_with_zero_21__16_  : 
                        (N55)? \xz.mem_with_zero_22__16_  : 
                        (N57)? \xz.mem_with_zero_23__16_  : 
                        (N59)? \xz.mem_with_zero_24__16_  : 
                        (N61)? \xz.mem_with_zero_25__16_  : 
                        (N63)? \xz.mem_with_zero_26__16_  : 
                        (N65)? \xz.mem_with_zero_27__16_  : 
                        (N67)? \xz.mem_with_zero_28__16_  : 
                        (N69)? \xz.mem_with_zero_29__16_  : 
                        (N71)? \xz.mem_with_zero_30__16_  : 
                        (N73)? \xz.mem_with_zero_31__16_  : 1'b0;
  assign r_data_o[15] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__15_  : 
                        (N46)? \xz.mem_with_zero_2__15_  : 
                        (N48)? \xz.mem_with_zero_3__15_  : 
                        (N50)? \xz.mem_with_zero_4__15_  : 
                        (N52)? \xz.mem_with_zero_5__15_  : 
                        (N54)? \xz.mem_with_zero_6__15_  : 
                        (N56)? \xz.mem_with_zero_7__15_  : 
                        (N58)? \xz.mem_with_zero_8__15_  : 
                        (N60)? \xz.mem_with_zero_9__15_  : 
                        (N62)? \xz.mem_with_zero_10__15_  : 
                        (N64)? \xz.mem_with_zero_11__15_  : 
                        (N66)? \xz.mem_with_zero_12__15_  : 
                        (N68)? \xz.mem_with_zero_13__15_  : 
                        (N70)? \xz.mem_with_zero_14__15_  : 
                        (N72)? \xz.mem_with_zero_15__15_  : 
                        (N43)? \xz.mem_with_zero_16__15_  : 
                        (N45)? \xz.mem_with_zero_17__15_  : 
                        (N47)? \xz.mem_with_zero_18__15_  : 
                        (N49)? \xz.mem_with_zero_19__15_  : 
                        (N51)? \xz.mem_with_zero_20__15_  : 
                        (N53)? \xz.mem_with_zero_21__15_  : 
                        (N55)? \xz.mem_with_zero_22__15_  : 
                        (N57)? \xz.mem_with_zero_23__15_  : 
                        (N59)? \xz.mem_with_zero_24__15_  : 
                        (N61)? \xz.mem_with_zero_25__15_  : 
                        (N63)? \xz.mem_with_zero_26__15_  : 
                        (N65)? \xz.mem_with_zero_27__15_  : 
                        (N67)? \xz.mem_with_zero_28__15_  : 
                        (N69)? \xz.mem_with_zero_29__15_  : 
                        (N71)? \xz.mem_with_zero_30__15_  : 
                        (N73)? \xz.mem_with_zero_31__15_  : 1'b0;
  assign r_data_o[14] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__14_  : 
                        (N46)? \xz.mem_with_zero_2__14_  : 
                        (N48)? \xz.mem_with_zero_3__14_  : 
                        (N50)? \xz.mem_with_zero_4__14_  : 
                        (N52)? \xz.mem_with_zero_5__14_  : 
                        (N54)? \xz.mem_with_zero_6__14_  : 
                        (N56)? \xz.mem_with_zero_7__14_  : 
                        (N58)? \xz.mem_with_zero_8__14_  : 
                        (N60)? \xz.mem_with_zero_9__14_  : 
                        (N62)? \xz.mem_with_zero_10__14_  : 
                        (N64)? \xz.mem_with_zero_11__14_  : 
                        (N66)? \xz.mem_with_zero_12__14_  : 
                        (N68)? \xz.mem_with_zero_13__14_  : 
                        (N70)? \xz.mem_with_zero_14__14_  : 
                        (N72)? \xz.mem_with_zero_15__14_  : 
                        (N43)? \xz.mem_with_zero_16__14_  : 
                        (N45)? \xz.mem_with_zero_17__14_  : 
                        (N47)? \xz.mem_with_zero_18__14_  : 
                        (N49)? \xz.mem_with_zero_19__14_  : 
                        (N51)? \xz.mem_with_zero_20__14_  : 
                        (N53)? \xz.mem_with_zero_21__14_  : 
                        (N55)? \xz.mem_with_zero_22__14_  : 
                        (N57)? \xz.mem_with_zero_23__14_  : 
                        (N59)? \xz.mem_with_zero_24__14_  : 
                        (N61)? \xz.mem_with_zero_25__14_  : 
                        (N63)? \xz.mem_with_zero_26__14_  : 
                        (N65)? \xz.mem_with_zero_27__14_  : 
                        (N67)? \xz.mem_with_zero_28__14_  : 
                        (N69)? \xz.mem_with_zero_29__14_  : 
                        (N71)? \xz.mem_with_zero_30__14_  : 
                        (N73)? \xz.mem_with_zero_31__14_  : 1'b0;
  assign r_data_o[13] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__13_  : 
                        (N46)? \xz.mem_with_zero_2__13_  : 
                        (N48)? \xz.mem_with_zero_3__13_  : 
                        (N50)? \xz.mem_with_zero_4__13_  : 
                        (N52)? \xz.mem_with_zero_5__13_  : 
                        (N54)? \xz.mem_with_zero_6__13_  : 
                        (N56)? \xz.mem_with_zero_7__13_  : 
                        (N58)? \xz.mem_with_zero_8__13_  : 
                        (N60)? \xz.mem_with_zero_9__13_  : 
                        (N62)? \xz.mem_with_zero_10__13_  : 
                        (N64)? \xz.mem_with_zero_11__13_  : 
                        (N66)? \xz.mem_with_zero_12__13_  : 
                        (N68)? \xz.mem_with_zero_13__13_  : 
                        (N70)? \xz.mem_with_zero_14__13_  : 
                        (N72)? \xz.mem_with_zero_15__13_  : 
                        (N43)? \xz.mem_with_zero_16__13_  : 
                        (N45)? \xz.mem_with_zero_17__13_  : 
                        (N47)? \xz.mem_with_zero_18__13_  : 
                        (N49)? \xz.mem_with_zero_19__13_  : 
                        (N51)? \xz.mem_with_zero_20__13_  : 
                        (N53)? \xz.mem_with_zero_21__13_  : 
                        (N55)? \xz.mem_with_zero_22__13_  : 
                        (N57)? \xz.mem_with_zero_23__13_  : 
                        (N59)? \xz.mem_with_zero_24__13_  : 
                        (N61)? \xz.mem_with_zero_25__13_  : 
                        (N63)? \xz.mem_with_zero_26__13_  : 
                        (N65)? \xz.mem_with_zero_27__13_  : 
                        (N67)? \xz.mem_with_zero_28__13_  : 
                        (N69)? \xz.mem_with_zero_29__13_  : 
                        (N71)? \xz.mem_with_zero_30__13_  : 
                        (N73)? \xz.mem_with_zero_31__13_  : 1'b0;
  assign r_data_o[12] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__12_  : 
                        (N46)? \xz.mem_with_zero_2__12_  : 
                        (N48)? \xz.mem_with_zero_3__12_  : 
                        (N50)? \xz.mem_with_zero_4__12_  : 
                        (N52)? \xz.mem_with_zero_5__12_  : 
                        (N54)? \xz.mem_with_zero_6__12_  : 
                        (N56)? \xz.mem_with_zero_7__12_  : 
                        (N58)? \xz.mem_with_zero_8__12_  : 
                        (N60)? \xz.mem_with_zero_9__12_  : 
                        (N62)? \xz.mem_with_zero_10__12_  : 
                        (N64)? \xz.mem_with_zero_11__12_  : 
                        (N66)? \xz.mem_with_zero_12__12_  : 
                        (N68)? \xz.mem_with_zero_13__12_  : 
                        (N70)? \xz.mem_with_zero_14__12_  : 
                        (N72)? \xz.mem_with_zero_15__12_  : 
                        (N43)? \xz.mem_with_zero_16__12_  : 
                        (N45)? \xz.mem_with_zero_17__12_  : 
                        (N47)? \xz.mem_with_zero_18__12_  : 
                        (N49)? \xz.mem_with_zero_19__12_  : 
                        (N51)? \xz.mem_with_zero_20__12_  : 
                        (N53)? \xz.mem_with_zero_21__12_  : 
                        (N55)? \xz.mem_with_zero_22__12_  : 
                        (N57)? \xz.mem_with_zero_23__12_  : 
                        (N59)? \xz.mem_with_zero_24__12_  : 
                        (N61)? \xz.mem_with_zero_25__12_  : 
                        (N63)? \xz.mem_with_zero_26__12_  : 
                        (N65)? \xz.mem_with_zero_27__12_  : 
                        (N67)? \xz.mem_with_zero_28__12_  : 
                        (N69)? \xz.mem_with_zero_29__12_  : 
                        (N71)? \xz.mem_with_zero_30__12_  : 
                        (N73)? \xz.mem_with_zero_31__12_  : 1'b0;
  assign r_data_o[11] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__11_  : 
                        (N46)? \xz.mem_with_zero_2__11_  : 
                        (N48)? \xz.mem_with_zero_3__11_  : 
                        (N50)? \xz.mem_with_zero_4__11_  : 
                        (N52)? \xz.mem_with_zero_5__11_  : 
                        (N54)? \xz.mem_with_zero_6__11_  : 
                        (N56)? \xz.mem_with_zero_7__11_  : 
                        (N58)? \xz.mem_with_zero_8__11_  : 
                        (N60)? \xz.mem_with_zero_9__11_  : 
                        (N62)? \xz.mem_with_zero_10__11_  : 
                        (N64)? \xz.mem_with_zero_11__11_  : 
                        (N66)? \xz.mem_with_zero_12__11_  : 
                        (N68)? \xz.mem_with_zero_13__11_  : 
                        (N70)? \xz.mem_with_zero_14__11_  : 
                        (N72)? \xz.mem_with_zero_15__11_  : 
                        (N43)? \xz.mem_with_zero_16__11_  : 
                        (N45)? \xz.mem_with_zero_17__11_  : 
                        (N47)? \xz.mem_with_zero_18__11_  : 
                        (N49)? \xz.mem_with_zero_19__11_  : 
                        (N51)? \xz.mem_with_zero_20__11_  : 
                        (N53)? \xz.mem_with_zero_21__11_  : 
                        (N55)? \xz.mem_with_zero_22__11_  : 
                        (N57)? \xz.mem_with_zero_23__11_  : 
                        (N59)? \xz.mem_with_zero_24__11_  : 
                        (N61)? \xz.mem_with_zero_25__11_  : 
                        (N63)? \xz.mem_with_zero_26__11_  : 
                        (N65)? \xz.mem_with_zero_27__11_  : 
                        (N67)? \xz.mem_with_zero_28__11_  : 
                        (N69)? \xz.mem_with_zero_29__11_  : 
                        (N71)? \xz.mem_with_zero_30__11_  : 
                        (N73)? \xz.mem_with_zero_31__11_  : 1'b0;
  assign r_data_o[10] = (N42)? 1'b0 : 
                        (N44)? \xz.mem_with_zero_1__10_  : 
                        (N46)? \xz.mem_with_zero_2__10_  : 
                        (N48)? \xz.mem_with_zero_3__10_  : 
                        (N50)? \xz.mem_with_zero_4__10_  : 
                        (N52)? \xz.mem_with_zero_5__10_  : 
                        (N54)? \xz.mem_with_zero_6__10_  : 
                        (N56)? \xz.mem_with_zero_7__10_  : 
                        (N58)? \xz.mem_with_zero_8__10_  : 
                        (N60)? \xz.mem_with_zero_9__10_  : 
                        (N62)? \xz.mem_with_zero_10__10_  : 
                        (N64)? \xz.mem_with_zero_11__10_  : 
                        (N66)? \xz.mem_with_zero_12__10_  : 
                        (N68)? \xz.mem_with_zero_13__10_  : 
                        (N70)? \xz.mem_with_zero_14__10_  : 
                        (N72)? \xz.mem_with_zero_15__10_  : 
                        (N43)? \xz.mem_with_zero_16__10_  : 
                        (N45)? \xz.mem_with_zero_17__10_  : 
                        (N47)? \xz.mem_with_zero_18__10_  : 
                        (N49)? \xz.mem_with_zero_19__10_  : 
                        (N51)? \xz.mem_with_zero_20__10_  : 
                        (N53)? \xz.mem_with_zero_21__10_  : 
                        (N55)? \xz.mem_with_zero_22__10_  : 
                        (N57)? \xz.mem_with_zero_23__10_  : 
                        (N59)? \xz.mem_with_zero_24__10_  : 
                        (N61)? \xz.mem_with_zero_25__10_  : 
                        (N63)? \xz.mem_with_zero_26__10_  : 
                        (N65)? \xz.mem_with_zero_27__10_  : 
                        (N67)? \xz.mem_with_zero_28__10_  : 
                        (N69)? \xz.mem_with_zero_29__10_  : 
                        (N71)? \xz.mem_with_zero_30__10_  : 
                        (N73)? \xz.mem_with_zero_31__10_  : 1'b0;
  assign r_data_o[9] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__9_  : 
                       (N46)? \xz.mem_with_zero_2__9_  : 
                       (N48)? \xz.mem_with_zero_3__9_  : 
                       (N50)? \xz.mem_with_zero_4__9_  : 
                       (N52)? \xz.mem_with_zero_5__9_  : 
                       (N54)? \xz.mem_with_zero_6__9_  : 
                       (N56)? \xz.mem_with_zero_7__9_  : 
                       (N58)? \xz.mem_with_zero_8__9_  : 
                       (N60)? \xz.mem_with_zero_9__9_  : 
                       (N62)? \xz.mem_with_zero_10__9_  : 
                       (N64)? \xz.mem_with_zero_11__9_  : 
                       (N66)? \xz.mem_with_zero_12__9_  : 
                       (N68)? \xz.mem_with_zero_13__9_  : 
                       (N70)? \xz.mem_with_zero_14__9_  : 
                       (N72)? \xz.mem_with_zero_15__9_  : 
                       (N43)? \xz.mem_with_zero_16__9_  : 
                       (N45)? \xz.mem_with_zero_17__9_  : 
                       (N47)? \xz.mem_with_zero_18__9_  : 
                       (N49)? \xz.mem_with_zero_19__9_  : 
                       (N51)? \xz.mem_with_zero_20__9_  : 
                       (N53)? \xz.mem_with_zero_21__9_  : 
                       (N55)? \xz.mem_with_zero_22__9_  : 
                       (N57)? \xz.mem_with_zero_23__9_  : 
                       (N59)? \xz.mem_with_zero_24__9_  : 
                       (N61)? \xz.mem_with_zero_25__9_  : 
                       (N63)? \xz.mem_with_zero_26__9_  : 
                       (N65)? \xz.mem_with_zero_27__9_  : 
                       (N67)? \xz.mem_with_zero_28__9_  : 
                       (N69)? \xz.mem_with_zero_29__9_  : 
                       (N71)? \xz.mem_with_zero_30__9_  : 
                       (N73)? \xz.mem_with_zero_31__9_  : 1'b0;
  assign r_data_o[8] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__8_  : 
                       (N46)? \xz.mem_with_zero_2__8_  : 
                       (N48)? \xz.mem_with_zero_3__8_  : 
                       (N50)? \xz.mem_with_zero_4__8_  : 
                       (N52)? \xz.mem_with_zero_5__8_  : 
                       (N54)? \xz.mem_with_zero_6__8_  : 
                       (N56)? \xz.mem_with_zero_7__8_  : 
                       (N58)? \xz.mem_with_zero_8__8_  : 
                       (N60)? \xz.mem_with_zero_9__8_  : 
                       (N62)? \xz.mem_with_zero_10__8_  : 
                       (N64)? \xz.mem_with_zero_11__8_  : 
                       (N66)? \xz.mem_with_zero_12__8_  : 
                       (N68)? \xz.mem_with_zero_13__8_  : 
                       (N70)? \xz.mem_with_zero_14__8_  : 
                       (N72)? \xz.mem_with_zero_15__8_  : 
                       (N43)? \xz.mem_with_zero_16__8_  : 
                       (N45)? \xz.mem_with_zero_17__8_  : 
                       (N47)? \xz.mem_with_zero_18__8_  : 
                       (N49)? \xz.mem_with_zero_19__8_  : 
                       (N51)? \xz.mem_with_zero_20__8_  : 
                       (N53)? \xz.mem_with_zero_21__8_  : 
                       (N55)? \xz.mem_with_zero_22__8_  : 
                       (N57)? \xz.mem_with_zero_23__8_  : 
                       (N59)? \xz.mem_with_zero_24__8_  : 
                       (N61)? \xz.mem_with_zero_25__8_  : 
                       (N63)? \xz.mem_with_zero_26__8_  : 
                       (N65)? \xz.mem_with_zero_27__8_  : 
                       (N67)? \xz.mem_with_zero_28__8_  : 
                       (N69)? \xz.mem_with_zero_29__8_  : 
                       (N71)? \xz.mem_with_zero_30__8_  : 
                       (N73)? \xz.mem_with_zero_31__8_  : 1'b0;
  assign r_data_o[7] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__7_  : 
                       (N46)? \xz.mem_with_zero_2__7_  : 
                       (N48)? \xz.mem_with_zero_3__7_  : 
                       (N50)? \xz.mem_with_zero_4__7_  : 
                       (N52)? \xz.mem_with_zero_5__7_  : 
                       (N54)? \xz.mem_with_zero_6__7_  : 
                       (N56)? \xz.mem_with_zero_7__7_  : 
                       (N58)? \xz.mem_with_zero_8__7_  : 
                       (N60)? \xz.mem_with_zero_9__7_  : 
                       (N62)? \xz.mem_with_zero_10__7_  : 
                       (N64)? \xz.mem_with_zero_11__7_  : 
                       (N66)? \xz.mem_with_zero_12__7_  : 
                       (N68)? \xz.mem_with_zero_13__7_  : 
                       (N70)? \xz.mem_with_zero_14__7_  : 
                       (N72)? \xz.mem_with_zero_15__7_  : 
                       (N43)? \xz.mem_with_zero_16__7_  : 
                       (N45)? \xz.mem_with_zero_17__7_  : 
                       (N47)? \xz.mem_with_zero_18__7_  : 
                       (N49)? \xz.mem_with_zero_19__7_  : 
                       (N51)? \xz.mem_with_zero_20__7_  : 
                       (N53)? \xz.mem_with_zero_21__7_  : 
                       (N55)? \xz.mem_with_zero_22__7_  : 
                       (N57)? \xz.mem_with_zero_23__7_  : 
                       (N59)? \xz.mem_with_zero_24__7_  : 
                       (N61)? \xz.mem_with_zero_25__7_  : 
                       (N63)? \xz.mem_with_zero_26__7_  : 
                       (N65)? \xz.mem_with_zero_27__7_  : 
                       (N67)? \xz.mem_with_zero_28__7_  : 
                       (N69)? \xz.mem_with_zero_29__7_  : 
                       (N71)? \xz.mem_with_zero_30__7_  : 
                       (N73)? \xz.mem_with_zero_31__7_  : 1'b0;
  assign r_data_o[6] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__6_  : 
                       (N46)? \xz.mem_with_zero_2__6_  : 
                       (N48)? \xz.mem_with_zero_3__6_  : 
                       (N50)? \xz.mem_with_zero_4__6_  : 
                       (N52)? \xz.mem_with_zero_5__6_  : 
                       (N54)? \xz.mem_with_zero_6__6_  : 
                       (N56)? \xz.mem_with_zero_7__6_  : 
                       (N58)? \xz.mem_with_zero_8__6_  : 
                       (N60)? \xz.mem_with_zero_9__6_  : 
                       (N62)? \xz.mem_with_zero_10__6_  : 
                       (N64)? \xz.mem_with_zero_11__6_  : 
                       (N66)? \xz.mem_with_zero_12__6_  : 
                       (N68)? \xz.mem_with_zero_13__6_  : 
                       (N70)? \xz.mem_with_zero_14__6_  : 
                       (N72)? \xz.mem_with_zero_15__6_  : 
                       (N43)? \xz.mem_with_zero_16__6_  : 
                       (N45)? \xz.mem_with_zero_17__6_  : 
                       (N47)? \xz.mem_with_zero_18__6_  : 
                       (N49)? \xz.mem_with_zero_19__6_  : 
                       (N51)? \xz.mem_with_zero_20__6_  : 
                       (N53)? \xz.mem_with_zero_21__6_  : 
                       (N55)? \xz.mem_with_zero_22__6_  : 
                       (N57)? \xz.mem_with_zero_23__6_  : 
                       (N59)? \xz.mem_with_zero_24__6_  : 
                       (N61)? \xz.mem_with_zero_25__6_  : 
                       (N63)? \xz.mem_with_zero_26__6_  : 
                       (N65)? \xz.mem_with_zero_27__6_  : 
                       (N67)? \xz.mem_with_zero_28__6_  : 
                       (N69)? \xz.mem_with_zero_29__6_  : 
                       (N71)? \xz.mem_with_zero_30__6_  : 
                       (N73)? \xz.mem_with_zero_31__6_  : 1'b0;
  assign r_data_o[5] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__5_  : 
                       (N46)? \xz.mem_with_zero_2__5_  : 
                       (N48)? \xz.mem_with_zero_3__5_  : 
                       (N50)? \xz.mem_with_zero_4__5_  : 
                       (N52)? \xz.mem_with_zero_5__5_  : 
                       (N54)? \xz.mem_with_zero_6__5_  : 
                       (N56)? \xz.mem_with_zero_7__5_  : 
                       (N58)? \xz.mem_with_zero_8__5_  : 
                       (N60)? \xz.mem_with_zero_9__5_  : 
                       (N62)? \xz.mem_with_zero_10__5_  : 
                       (N64)? \xz.mem_with_zero_11__5_  : 
                       (N66)? \xz.mem_with_zero_12__5_  : 
                       (N68)? \xz.mem_with_zero_13__5_  : 
                       (N70)? \xz.mem_with_zero_14__5_  : 
                       (N72)? \xz.mem_with_zero_15__5_  : 
                       (N43)? \xz.mem_with_zero_16__5_  : 
                       (N45)? \xz.mem_with_zero_17__5_  : 
                       (N47)? \xz.mem_with_zero_18__5_  : 
                       (N49)? \xz.mem_with_zero_19__5_  : 
                       (N51)? \xz.mem_with_zero_20__5_  : 
                       (N53)? \xz.mem_with_zero_21__5_  : 
                       (N55)? \xz.mem_with_zero_22__5_  : 
                       (N57)? \xz.mem_with_zero_23__5_  : 
                       (N59)? \xz.mem_with_zero_24__5_  : 
                       (N61)? \xz.mem_with_zero_25__5_  : 
                       (N63)? \xz.mem_with_zero_26__5_  : 
                       (N65)? \xz.mem_with_zero_27__5_  : 
                       (N67)? \xz.mem_with_zero_28__5_  : 
                       (N69)? \xz.mem_with_zero_29__5_  : 
                       (N71)? \xz.mem_with_zero_30__5_  : 
                       (N73)? \xz.mem_with_zero_31__5_  : 1'b0;
  assign r_data_o[4] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__4_  : 
                       (N46)? \xz.mem_with_zero_2__4_  : 
                       (N48)? \xz.mem_with_zero_3__4_  : 
                       (N50)? \xz.mem_with_zero_4__4_  : 
                       (N52)? \xz.mem_with_zero_5__4_  : 
                       (N54)? \xz.mem_with_zero_6__4_  : 
                       (N56)? \xz.mem_with_zero_7__4_  : 
                       (N58)? \xz.mem_with_zero_8__4_  : 
                       (N60)? \xz.mem_with_zero_9__4_  : 
                       (N62)? \xz.mem_with_zero_10__4_  : 
                       (N64)? \xz.mem_with_zero_11__4_  : 
                       (N66)? \xz.mem_with_zero_12__4_  : 
                       (N68)? \xz.mem_with_zero_13__4_  : 
                       (N70)? \xz.mem_with_zero_14__4_  : 
                       (N72)? \xz.mem_with_zero_15__4_  : 
                       (N43)? \xz.mem_with_zero_16__4_  : 
                       (N45)? \xz.mem_with_zero_17__4_  : 
                       (N47)? \xz.mem_with_zero_18__4_  : 
                       (N49)? \xz.mem_with_zero_19__4_  : 
                       (N51)? \xz.mem_with_zero_20__4_  : 
                       (N53)? \xz.mem_with_zero_21__4_  : 
                       (N55)? \xz.mem_with_zero_22__4_  : 
                       (N57)? \xz.mem_with_zero_23__4_  : 
                       (N59)? \xz.mem_with_zero_24__4_  : 
                       (N61)? \xz.mem_with_zero_25__4_  : 
                       (N63)? \xz.mem_with_zero_26__4_  : 
                       (N65)? \xz.mem_with_zero_27__4_  : 
                       (N67)? \xz.mem_with_zero_28__4_  : 
                       (N69)? \xz.mem_with_zero_29__4_  : 
                       (N71)? \xz.mem_with_zero_30__4_  : 
                       (N73)? \xz.mem_with_zero_31__4_  : 1'b0;
  assign r_data_o[3] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__3_  : 
                       (N46)? \xz.mem_with_zero_2__3_  : 
                       (N48)? \xz.mem_with_zero_3__3_  : 
                       (N50)? \xz.mem_with_zero_4__3_  : 
                       (N52)? \xz.mem_with_zero_5__3_  : 
                       (N54)? \xz.mem_with_zero_6__3_  : 
                       (N56)? \xz.mem_with_zero_7__3_  : 
                       (N58)? \xz.mem_with_zero_8__3_  : 
                       (N60)? \xz.mem_with_zero_9__3_  : 
                       (N62)? \xz.mem_with_zero_10__3_  : 
                       (N64)? \xz.mem_with_zero_11__3_  : 
                       (N66)? \xz.mem_with_zero_12__3_  : 
                       (N68)? \xz.mem_with_zero_13__3_  : 
                       (N70)? \xz.mem_with_zero_14__3_  : 
                       (N72)? \xz.mem_with_zero_15__3_  : 
                       (N43)? \xz.mem_with_zero_16__3_  : 
                       (N45)? \xz.mem_with_zero_17__3_  : 
                       (N47)? \xz.mem_with_zero_18__3_  : 
                       (N49)? \xz.mem_with_zero_19__3_  : 
                       (N51)? \xz.mem_with_zero_20__3_  : 
                       (N53)? \xz.mem_with_zero_21__3_  : 
                       (N55)? \xz.mem_with_zero_22__3_  : 
                       (N57)? \xz.mem_with_zero_23__3_  : 
                       (N59)? \xz.mem_with_zero_24__3_  : 
                       (N61)? \xz.mem_with_zero_25__3_  : 
                       (N63)? \xz.mem_with_zero_26__3_  : 
                       (N65)? \xz.mem_with_zero_27__3_  : 
                       (N67)? \xz.mem_with_zero_28__3_  : 
                       (N69)? \xz.mem_with_zero_29__3_  : 
                       (N71)? \xz.mem_with_zero_30__3_  : 
                       (N73)? \xz.mem_with_zero_31__3_  : 1'b0;
  assign r_data_o[2] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__2_  : 
                       (N46)? \xz.mem_with_zero_2__2_  : 
                       (N48)? \xz.mem_with_zero_3__2_  : 
                       (N50)? \xz.mem_with_zero_4__2_  : 
                       (N52)? \xz.mem_with_zero_5__2_  : 
                       (N54)? \xz.mem_with_zero_6__2_  : 
                       (N56)? \xz.mem_with_zero_7__2_  : 
                       (N58)? \xz.mem_with_zero_8__2_  : 
                       (N60)? \xz.mem_with_zero_9__2_  : 
                       (N62)? \xz.mem_with_zero_10__2_  : 
                       (N64)? \xz.mem_with_zero_11__2_  : 
                       (N66)? \xz.mem_with_zero_12__2_  : 
                       (N68)? \xz.mem_with_zero_13__2_  : 
                       (N70)? \xz.mem_with_zero_14__2_  : 
                       (N72)? \xz.mem_with_zero_15__2_  : 
                       (N43)? \xz.mem_with_zero_16__2_  : 
                       (N45)? \xz.mem_with_zero_17__2_  : 
                       (N47)? \xz.mem_with_zero_18__2_  : 
                       (N49)? \xz.mem_with_zero_19__2_  : 
                       (N51)? \xz.mem_with_zero_20__2_  : 
                       (N53)? \xz.mem_with_zero_21__2_  : 
                       (N55)? \xz.mem_with_zero_22__2_  : 
                       (N57)? \xz.mem_with_zero_23__2_  : 
                       (N59)? \xz.mem_with_zero_24__2_  : 
                       (N61)? \xz.mem_with_zero_25__2_  : 
                       (N63)? \xz.mem_with_zero_26__2_  : 
                       (N65)? \xz.mem_with_zero_27__2_  : 
                       (N67)? \xz.mem_with_zero_28__2_  : 
                       (N69)? \xz.mem_with_zero_29__2_  : 
                       (N71)? \xz.mem_with_zero_30__2_  : 
                       (N73)? \xz.mem_with_zero_31__2_  : 1'b0;
  assign r_data_o[1] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__1_  : 
                       (N46)? \xz.mem_with_zero_2__1_  : 
                       (N48)? \xz.mem_with_zero_3__1_  : 
                       (N50)? \xz.mem_with_zero_4__1_  : 
                       (N52)? \xz.mem_with_zero_5__1_  : 
                       (N54)? \xz.mem_with_zero_6__1_  : 
                       (N56)? \xz.mem_with_zero_7__1_  : 
                       (N58)? \xz.mem_with_zero_8__1_  : 
                       (N60)? \xz.mem_with_zero_9__1_  : 
                       (N62)? \xz.mem_with_zero_10__1_  : 
                       (N64)? \xz.mem_with_zero_11__1_  : 
                       (N66)? \xz.mem_with_zero_12__1_  : 
                       (N68)? \xz.mem_with_zero_13__1_  : 
                       (N70)? \xz.mem_with_zero_14__1_  : 
                       (N72)? \xz.mem_with_zero_15__1_  : 
                       (N43)? \xz.mem_with_zero_16__1_  : 
                       (N45)? \xz.mem_with_zero_17__1_  : 
                       (N47)? \xz.mem_with_zero_18__1_  : 
                       (N49)? \xz.mem_with_zero_19__1_  : 
                       (N51)? \xz.mem_with_zero_20__1_  : 
                       (N53)? \xz.mem_with_zero_21__1_  : 
                       (N55)? \xz.mem_with_zero_22__1_  : 
                       (N57)? \xz.mem_with_zero_23__1_  : 
                       (N59)? \xz.mem_with_zero_24__1_  : 
                       (N61)? \xz.mem_with_zero_25__1_  : 
                       (N63)? \xz.mem_with_zero_26__1_  : 
                       (N65)? \xz.mem_with_zero_27__1_  : 
                       (N67)? \xz.mem_with_zero_28__1_  : 
                       (N69)? \xz.mem_with_zero_29__1_  : 
                       (N71)? \xz.mem_with_zero_30__1_  : 
                       (N73)? \xz.mem_with_zero_31__1_  : 1'b0;
  assign r_data_o[0] = (N42)? 1'b0 : 
                       (N44)? \xz.mem_with_zero_1__0_  : 
                       (N46)? \xz.mem_with_zero_2__0_  : 
                       (N48)? \xz.mem_with_zero_3__0_  : 
                       (N50)? \xz.mem_with_zero_4__0_  : 
                       (N52)? \xz.mem_with_zero_5__0_  : 
                       (N54)? \xz.mem_with_zero_6__0_  : 
                       (N56)? \xz.mem_with_zero_7__0_  : 
                       (N58)? \xz.mem_with_zero_8__0_  : 
                       (N60)? \xz.mem_with_zero_9__0_  : 
                       (N62)? \xz.mem_with_zero_10__0_  : 
                       (N64)? \xz.mem_with_zero_11__0_  : 
                       (N66)? \xz.mem_with_zero_12__0_  : 
                       (N68)? \xz.mem_with_zero_13__0_  : 
                       (N70)? \xz.mem_with_zero_14__0_  : 
                       (N72)? \xz.mem_with_zero_15__0_  : 
                       (N43)? \xz.mem_with_zero_16__0_  : 
                       (N45)? \xz.mem_with_zero_17__0_  : 
                       (N47)? \xz.mem_with_zero_18__0_  : 
                       (N49)? \xz.mem_with_zero_19__0_  : 
                       (N51)? \xz.mem_with_zero_20__0_  : 
                       (N53)? \xz.mem_with_zero_21__0_  : 
                       (N55)? \xz.mem_with_zero_22__0_  : 
                       (N57)? \xz.mem_with_zero_23__0_  : 
                       (N59)? \xz.mem_with_zero_24__0_  : 
                       (N61)? \xz.mem_with_zero_25__0_  : 
                       (N63)? \xz.mem_with_zero_26__0_  : 
                       (N65)? \xz.mem_with_zero_27__0_  : 
                       (N67)? \xz.mem_with_zero_28__0_  : 
                       (N69)? \xz.mem_with_zero_29__0_  : 
                       (N71)? \xz.mem_with_zero_30__0_  : 
                       (N73)? \xz.mem_with_zero_31__0_  : 1'b0;
  assign r_data_o[63] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__31_  : 
                        (N111)? \xz.mem_with_zero_2__31_  : 
                        (N113)? \xz.mem_with_zero_3__31_  : 
                        (N115)? \xz.mem_with_zero_4__31_  : 
                        (N117)? \xz.mem_with_zero_5__31_  : 
                        (N119)? \xz.mem_with_zero_6__31_  : 
                        (N121)? \xz.mem_with_zero_7__31_  : 
                        (N123)? \xz.mem_with_zero_8__31_  : 
                        (N125)? \xz.mem_with_zero_9__31_  : 
                        (N127)? \xz.mem_with_zero_10__31_  : 
                        (N129)? \xz.mem_with_zero_11__31_  : 
                        (N131)? \xz.mem_with_zero_12__31_  : 
                        (N133)? \xz.mem_with_zero_13__31_  : 
                        (N135)? \xz.mem_with_zero_14__31_  : 
                        (N137)? \xz.mem_with_zero_15__31_  : 
                        (N108)? \xz.mem_with_zero_16__31_  : 
                        (N110)? \xz.mem_with_zero_17__31_  : 
                        (N112)? \xz.mem_with_zero_18__31_  : 
                        (N114)? \xz.mem_with_zero_19__31_  : 
                        (N116)? \xz.mem_with_zero_20__31_  : 
                        (N118)? \xz.mem_with_zero_21__31_  : 
                        (N120)? \xz.mem_with_zero_22__31_  : 
                        (N122)? \xz.mem_with_zero_23__31_  : 
                        (N124)? \xz.mem_with_zero_24__31_  : 
                        (N126)? \xz.mem_with_zero_25__31_  : 
                        (N128)? \xz.mem_with_zero_26__31_  : 
                        (N130)? \xz.mem_with_zero_27__31_  : 
                        (N132)? \xz.mem_with_zero_28__31_  : 
                        (N134)? \xz.mem_with_zero_29__31_  : 
                        (N136)? \xz.mem_with_zero_30__31_  : 
                        (N138)? \xz.mem_with_zero_31__31_  : 1'b0;
  assign r_data_o[62] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__30_  : 
                        (N111)? \xz.mem_with_zero_2__30_  : 
                        (N113)? \xz.mem_with_zero_3__30_  : 
                        (N115)? \xz.mem_with_zero_4__30_  : 
                        (N117)? \xz.mem_with_zero_5__30_  : 
                        (N119)? \xz.mem_with_zero_6__30_  : 
                        (N121)? \xz.mem_with_zero_7__30_  : 
                        (N123)? \xz.mem_with_zero_8__30_  : 
                        (N125)? \xz.mem_with_zero_9__30_  : 
                        (N127)? \xz.mem_with_zero_10__30_  : 
                        (N129)? \xz.mem_with_zero_11__30_  : 
                        (N131)? \xz.mem_with_zero_12__30_  : 
                        (N133)? \xz.mem_with_zero_13__30_  : 
                        (N135)? \xz.mem_with_zero_14__30_  : 
                        (N137)? \xz.mem_with_zero_15__30_  : 
                        (N108)? \xz.mem_with_zero_16__30_  : 
                        (N110)? \xz.mem_with_zero_17__30_  : 
                        (N112)? \xz.mem_with_zero_18__30_  : 
                        (N114)? \xz.mem_with_zero_19__30_  : 
                        (N116)? \xz.mem_with_zero_20__30_  : 
                        (N118)? \xz.mem_with_zero_21__30_  : 
                        (N120)? \xz.mem_with_zero_22__30_  : 
                        (N122)? \xz.mem_with_zero_23__30_  : 
                        (N124)? \xz.mem_with_zero_24__30_  : 
                        (N126)? \xz.mem_with_zero_25__30_  : 
                        (N128)? \xz.mem_with_zero_26__30_  : 
                        (N130)? \xz.mem_with_zero_27__30_  : 
                        (N132)? \xz.mem_with_zero_28__30_  : 
                        (N134)? \xz.mem_with_zero_29__30_  : 
                        (N136)? \xz.mem_with_zero_30__30_  : 
                        (N138)? \xz.mem_with_zero_31__30_  : 1'b0;
  assign r_data_o[61] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__29_  : 
                        (N111)? \xz.mem_with_zero_2__29_  : 
                        (N113)? \xz.mem_with_zero_3__29_  : 
                        (N115)? \xz.mem_with_zero_4__29_  : 
                        (N117)? \xz.mem_with_zero_5__29_  : 
                        (N119)? \xz.mem_with_zero_6__29_  : 
                        (N121)? \xz.mem_with_zero_7__29_  : 
                        (N123)? \xz.mem_with_zero_8__29_  : 
                        (N125)? \xz.mem_with_zero_9__29_  : 
                        (N127)? \xz.mem_with_zero_10__29_  : 
                        (N129)? \xz.mem_with_zero_11__29_  : 
                        (N131)? \xz.mem_with_zero_12__29_  : 
                        (N133)? \xz.mem_with_zero_13__29_  : 
                        (N135)? \xz.mem_with_zero_14__29_  : 
                        (N137)? \xz.mem_with_zero_15__29_  : 
                        (N108)? \xz.mem_with_zero_16__29_  : 
                        (N110)? \xz.mem_with_zero_17__29_  : 
                        (N112)? \xz.mem_with_zero_18__29_  : 
                        (N114)? \xz.mem_with_zero_19__29_  : 
                        (N116)? \xz.mem_with_zero_20__29_  : 
                        (N118)? \xz.mem_with_zero_21__29_  : 
                        (N120)? \xz.mem_with_zero_22__29_  : 
                        (N122)? \xz.mem_with_zero_23__29_  : 
                        (N124)? \xz.mem_with_zero_24__29_  : 
                        (N126)? \xz.mem_with_zero_25__29_  : 
                        (N128)? \xz.mem_with_zero_26__29_  : 
                        (N130)? \xz.mem_with_zero_27__29_  : 
                        (N132)? \xz.mem_with_zero_28__29_  : 
                        (N134)? \xz.mem_with_zero_29__29_  : 
                        (N136)? \xz.mem_with_zero_30__29_  : 
                        (N138)? \xz.mem_with_zero_31__29_  : 1'b0;
  assign r_data_o[60] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__28_  : 
                        (N111)? \xz.mem_with_zero_2__28_  : 
                        (N113)? \xz.mem_with_zero_3__28_  : 
                        (N115)? \xz.mem_with_zero_4__28_  : 
                        (N117)? \xz.mem_with_zero_5__28_  : 
                        (N119)? \xz.mem_with_zero_6__28_  : 
                        (N121)? \xz.mem_with_zero_7__28_  : 
                        (N123)? \xz.mem_with_zero_8__28_  : 
                        (N125)? \xz.mem_with_zero_9__28_  : 
                        (N127)? \xz.mem_with_zero_10__28_  : 
                        (N129)? \xz.mem_with_zero_11__28_  : 
                        (N131)? \xz.mem_with_zero_12__28_  : 
                        (N133)? \xz.mem_with_zero_13__28_  : 
                        (N135)? \xz.mem_with_zero_14__28_  : 
                        (N137)? \xz.mem_with_zero_15__28_  : 
                        (N108)? \xz.mem_with_zero_16__28_  : 
                        (N110)? \xz.mem_with_zero_17__28_  : 
                        (N112)? \xz.mem_with_zero_18__28_  : 
                        (N114)? \xz.mem_with_zero_19__28_  : 
                        (N116)? \xz.mem_with_zero_20__28_  : 
                        (N118)? \xz.mem_with_zero_21__28_  : 
                        (N120)? \xz.mem_with_zero_22__28_  : 
                        (N122)? \xz.mem_with_zero_23__28_  : 
                        (N124)? \xz.mem_with_zero_24__28_  : 
                        (N126)? \xz.mem_with_zero_25__28_  : 
                        (N128)? \xz.mem_with_zero_26__28_  : 
                        (N130)? \xz.mem_with_zero_27__28_  : 
                        (N132)? \xz.mem_with_zero_28__28_  : 
                        (N134)? \xz.mem_with_zero_29__28_  : 
                        (N136)? \xz.mem_with_zero_30__28_  : 
                        (N138)? \xz.mem_with_zero_31__28_  : 1'b0;
  assign r_data_o[59] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__27_  : 
                        (N111)? \xz.mem_with_zero_2__27_  : 
                        (N113)? \xz.mem_with_zero_3__27_  : 
                        (N115)? \xz.mem_with_zero_4__27_  : 
                        (N117)? \xz.mem_with_zero_5__27_  : 
                        (N119)? \xz.mem_with_zero_6__27_  : 
                        (N121)? \xz.mem_with_zero_7__27_  : 
                        (N123)? \xz.mem_with_zero_8__27_  : 
                        (N125)? \xz.mem_with_zero_9__27_  : 
                        (N127)? \xz.mem_with_zero_10__27_  : 
                        (N129)? \xz.mem_with_zero_11__27_  : 
                        (N131)? \xz.mem_with_zero_12__27_  : 
                        (N133)? \xz.mem_with_zero_13__27_  : 
                        (N135)? \xz.mem_with_zero_14__27_  : 
                        (N137)? \xz.mem_with_zero_15__27_  : 
                        (N108)? \xz.mem_with_zero_16__27_  : 
                        (N110)? \xz.mem_with_zero_17__27_  : 
                        (N112)? \xz.mem_with_zero_18__27_  : 
                        (N114)? \xz.mem_with_zero_19__27_  : 
                        (N116)? \xz.mem_with_zero_20__27_  : 
                        (N118)? \xz.mem_with_zero_21__27_  : 
                        (N120)? \xz.mem_with_zero_22__27_  : 
                        (N122)? \xz.mem_with_zero_23__27_  : 
                        (N124)? \xz.mem_with_zero_24__27_  : 
                        (N126)? \xz.mem_with_zero_25__27_  : 
                        (N128)? \xz.mem_with_zero_26__27_  : 
                        (N130)? \xz.mem_with_zero_27__27_  : 
                        (N132)? \xz.mem_with_zero_28__27_  : 
                        (N134)? \xz.mem_with_zero_29__27_  : 
                        (N136)? \xz.mem_with_zero_30__27_  : 
                        (N138)? \xz.mem_with_zero_31__27_  : 1'b0;
  assign r_data_o[58] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__26_  : 
                        (N111)? \xz.mem_with_zero_2__26_  : 
                        (N113)? \xz.mem_with_zero_3__26_  : 
                        (N115)? \xz.mem_with_zero_4__26_  : 
                        (N117)? \xz.mem_with_zero_5__26_  : 
                        (N119)? \xz.mem_with_zero_6__26_  : 
                        (N121)? \xz.mem_with_zero_7__26_  : 
                        (N123)? \xz.mem_with_zero_8__26_  : 
                        (N125)? \xz.mem_with_zero_9__26_  : 
                        (N127)? \xz.mem_with_zero_10__26_  : 
                        (N129)? \xz.mem_with_zero_11__26_  : 
                        (N131)? \xz.mem_with_zero_12__26_  : 
                        (N133)? \xz.mem_with_zero_13__26_  : 
                        (N135)? \xz.mem_with_zero_14__26_  : 
                        (N137)? \xz.mem_with_zero_15__26_  : 
                        (N108)? \xz.mem_with_zero_16__26_  : 
                        (N110)? \xz.mem_with_zero_17__26_  : 
                        (N112)? \xz.mem_with_zero_18__26_  : 
                        (N114)? \xz.mem_with_zero_19__26_  : 
                        (N116)? \xz.mem_with_zero_20__26_  : 
                        (N118)? \xz.mem_with_zero_21__26_  : 
                        (N120)? \xz.mem_with_zero_22__26_  : 
                        (N122)? \xz.mem_with_zero_23__26_  : 
                        (N124)? \xz.mem_with_zero_24__26_  : 
                        (N126)? \xz.mem_with_zero_25__26_  : 
                        (N128)? \xz.mem_with_zero_26__26_  : 
                        (N130)? \xz.mem_with_zero_27__26_  : 
                        (N132)? \xz.mem_with_zero_28__26_  : 
                        (N134)? \xz.mem_with_zero_29__26_  : 
                        (N136)? \xz.mem_with_zero_30__26_  : 
                        (N138)? \xz.mem_with_zero_31__26_  : 1'b0;
  assign r_data_o[57] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__25_  : 
                        (N111)? \xz.mem_with_zero_2__25_  : 
                        (N113)? \xz.mem_with_zero_3__25_  : 
                        (N115)? \xz.mem_with_zero_4__25_  : 
                        (N117)? \xz.mem_with_zero_5__25_  : 
                        (N119)? \xz.mem_with_zero_6__25_  : 
                        (N121)? \xz.mem_with_zero_7__25_  : 
                        (N123)? \xz.mem_with_zero_8__25_  : 
                        (N125)? \xz.mem_with_zero_9__25_  : 
                        (N127)? \xz.mem_with_zero_10__25_  : 
                        (N129)? \xz.mem_with_zero_11__25_  : 
                        (N131)? \xz.mem_with_zero_12__25_  : 
                        (N133)? \xz.mem_with_zero_13__25_  : 
                        (N135)? \xz.mem_with_zero_14__25_  : 
                        (N137)? \xz.mem_with_zero_15__25_  : 
                        (N108)? \xz.mem_with_zero_16__25_  : 
                        (N110)? \xz.mem_with_zero_17__25_  : 
                        (N112)? \xz.mem_with_zero_18__25_  : 
                        (N114)? \xz.mem_with_zero_19__25_  : 
                        (N116)? \xz.mem_with_zero_20__25_  : 
                        (N118)? \xz.mem_with_zero_21__25_  : 
                        (N120)? \xz.mem_with_zero_22__25_  : 
                        (N122)? \xz.mem_with_zero_23__25_  : 
                        (N124)? \xz.mem_with_zero_24__25_  : 
                        (N126)? \xz.mem_with_zero_25__25_  : 
                        (N128)? \xz.mem_with_zero_26__25_  : 
                        (N130)? \xz.mem_with_zero_27__25_  : 
                        (N132)? \xz.mem_with_zero_28__25_  : 
                        (N134)? \xz.mem_with_zero_29__25_  : 
                        (N136)? \xz.mem_with_zero_30__25_  : 
                        (N138)? \xz.mem_with_zero_31__25_  : 1'b0;
  assign r_data_o[56] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__24_  : 
                        (N111)? \xz.mem_with_zero_2__24_  : 
                        (N113)? \xz.mem_with_zero_3__24_  : 
                        (N115)? \xz.mem_with_zero_4__24_  : 
                        (N117)? \xz.mem_with_zero_5__24_  : 
                        (N119)? \xz.mem_with_zero_6__24_  : 
                        (N121)? \xz.mem_with_zero_7__24_  : 
                        (N123)? \xz.mem_with_zero_8__24_  : 
                        (N125)? \xz.mem_with_zero_9__24_  : 
                        (N127)? \xz.mem_with_zero_10__24_  : 
                        (N129)? \xz.mem_with_zero_11__24_  : 
                        (N131)? \xz.mem_with_zero_12__24_  : 
                        (N133)? \xz.mem_with_zero_13__24_  : 
                        (N135)? \xz.mem_with_zero_14__24_  : 
                        (N137)? \xz.mem_with_zero_15__24_  : 
                        (N108)? \xz.mem_with_zero_16__24_  : 
                        (N110)? \xz.mem_with_zero_17__24_  : 
                        (N112)? \xz.mem_with_zero_18__24_  : 
                        (N114)? \xz.mem_with_zero_19__24_  : 
                        (N116)? \xz.mem_with_zero_20__24_  : 
                        (N118)? \xz.mem_with_zero_21__24_  : 
                        (N120)? \xz.mem_with_zero_22__24_  : 
                        (N122)? \xz.mem_with_zero_23__24_  : 
                        (N124)? \xz.mem_with_zero_24__24_  : 
                        (N126)? \xz.mem_with_zero_25__24_  : 
                        (N128)? \xz.mem_with_zero_26__24_  : 
                        (N130)? \xz.mem_with_zero_27__24_  : 
                        (N132)? \xz.mem_with_zero_28__24_  : 
                        (N134)? \xz.mem_with_zero_29__24_  : 
                        (N136)? \xz.mem_with_zero_30__24_  : 
                        (N138)? \xz.mem_with_zero_31__24_  : 1'b0;
  assign r_data_o[55] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__23_  : 
                        (N111)? \xz.mem_with_zero_2__23_  : 
                        (N113)? \xz.mem_with_zero_3__23_  : 
                        (N115)? \xz.mem_with_zero_4__23_  : 
                        (N117)? \xz.mem_with_zero_5__23_  : 
                        (N119)? \xz.mem_with_zero_6__23_  : 
                        (N121)? \xz.mem_with_zero_7__23_  : 
                        (N123)? \xz.mem_with_zero_8__23_  : 
                        (N125)? \xz.mem_with_zero_9__23_  : 
                        (N127)? \xz.mem_with_zero_10__23_  : 
                        (N129)? \xz.mem_with_zero_11__23_  : 
                        (N131)? \xz.mem_with_zero_12__23_  : 
                        (N133)? \xz.mem_with_zero_13__23_  : 
                        (N135)? \xz.mem_with_zero_14__23_  : 
                        (N137)? \xz.mem_with_zero_15__23_  : 
                        (N108)? \xz.mem_with_zero_16__23_  : 
                        (N110)? \xz.mem_with_zero_17__23_  : 
                        (N112)? \xz.mem_with_zero_18__23_  : 
                        (N114)? \xz.mem_with_zero_19__23_  : 
                        (N116)? \xz.mem_with_zero_20__23_  : 
                        (N118)? \xz.mem_with_zero_21__23_  : 
                        (N120)? \xz.mem_with_zero_22__23_  : 
                        (N122)? \xz.mem_with_zero_23__23_  : 
                        (N124)? \xz.mem_with_zero_24__23_  : 
                        (N126)? \xz.mem_with_zero_25__23_  : 
                        (N128)? \xz.mem_with_zero_26__23_  : 
                        (N130)? \xz.mem_with_zero_27__23_  : 
                        (N132)? \xz.mem_with_zero_28__23_  : 
                        (N134)? \xz.mem_with_zero_29__23_  : 
                        (N136)? \xz.mem_with_zero_30__23_  : 
                        (N138)? \xz.mem_with_zero_31__23_  : 1'b0;
  assign r_data_o[54] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__22_  : 
                        (N111)? \xz.mem_with_zero_2__22_  : 
                        (N113)? \xz.mem_with_zero_3__22_  : 
                        (N115)? \xz.mem_with_zero_4__22_  : 
                        (N117)? \xz.mem_with_zero_5__22_  : 
                        (N119)? \xz.mem_with_zero_6__22_  : 
                        (N121)? \xz.mem_with_zero_7__22_  : 
                        (N123)? \xz.mem_with_zero_8__22_  : 
                        (N125)? \xz.mem_with_zero_9__22_  : 
                        (N127)? \xz.mem_with_zero_10__22_  : 
                        (N129)? \xz.mem_with_zero_11__22_  : 
                        (N131)? \xz.mem_with_zero_12__22_  : 
                        (N133)? \xz.mem_with_zero_13__22_  : 
                        (N135)? \xz.mem_with_zero_14__22_  : 
                        (N137)? \xz.mem_with_zero_15__22_  : 
                        (N108)? \xz.mem_with_zero_16__22_  : 
                        (N110)? \xz.mem_with_zero_17__22_  : 
                        (N112)? \xz.mem_with_zero_18__22_  : 
                        (N114)? \xz.mem_with_zero_19__22_  : 
                        (N116)? \xz.mem_with_zero_20__22_  : 
                        (N118)? \xz.mem_with_zero_21__22_  : 
                        (N120)? \xz.mem_with_zero_22__22_  : 
                        (N122)? \xz.mem_with_zero_23__22_  : 
                        (N124)? \xz.mem_with_zero_24__22_  : 
                        (N126)? \xz.mem_with_zero_25__22_  : 
                        (N128)? \xz.mem_with_zero_26__22_  : 
                        (N130)? \xz.mem_with_zero_27__22_  : 
                        (N132)? \xz.mem_with_zero_28__22_  : 
                        (N134)? \xz.mem_with_zero_29__22_  : 
                        (N136)? \xz.mem_with_zero_30__22_  : 
                        (N138)? \xz.mem_with_zero_31__22_  : 1'b0;
  assign r_data_o[53] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__21_  : 
                        (N111)? \xz.mem_with_zero_2__21_  : 
                        (N113)? \xz.mem_with_zero_3__21_  : 
                        (N115)? \xz.mem_with_zero_4__21_  : 
                        (N117)? \xz.mem_with_zero_5__21_  : 
                        (N119)? \xz.mem_with_zero_6__21_  : 
                        (N121)? \xz.mem_with_zero_7__21_  : 
                        (N123)? \xz.mem_with_zero_8__21_  : 
                        (N125)? \xz.mem_with_zero_9__21_  : 
                        (N127)? \xz.mem_with_zero_10__21_  : 
                        (N129)? \xz.mem_with_zero_11__21_  : 
                        (N131)? \xz.mem_with_zero_12__21_  : 
                        (N133)? \xz.mem_with_zero_13__21_  : 
                        (N135)? \xz.mem_with_zero_14__21_  : 
                        (N137)? \xz.mem_with_zero_15__21_  : 
                        (N108)? \xz.mem_with_zero_16__21_  : 
                        (N110)? \xz.mem_with_zero_17__21_  : 
                        (N112)? \xz.mem_with_zero_18__21_  : 
                        (N114)? \xz.mem_with_zero_19__21_  : 
                        (N116)? \xz.mem_with_zero_20__21_  : 
                        (N118)? \xz.mem_with_zero_21__21_  : 
                        (N120)? \xz.mem_with_zero_22__21_  : 
                        (N122)? \xz.mem_with_zero_23__21_  : 
                        (N124)? \xz.mem_with_zero_24__21_  : 
                        (N126)? \xz.mem_with_zero_25__21_  : 
                        (N128)? \xz.mem_with_zero_26__21_  : 
                        (N130)? \xz.mem_with_zero_27__21_  : 
                        (N132)? \xz.mem_with_zero_28__21_  : 
                        (N134)? \xz.mem_with_zero_29__21_  : 
                        (N136)? \xz.mem_with_zero_30__21_  : 
                        (N138)? \xz.mem_with_zero_31__21_  : 1'b0;
  assign r_data_o[52] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__20_  : 
                        (N111)? \xz.mem_with_zero_2__20_  : 
                        (N113)? \xz.mem_with_zero_3__20_  : 
                        (N115)? \xz.mem_with_zero_4__20_  : 
                        (N117)? \xz.mem_with_zero_5__20_  : 
                        (N119)? \xz.mem_with_zero_6__20_  : 
                        (N121)? \xz.mem_with_zero_7__20_  : 
                        (N123)? \xz.mem_with_zero_8__20_  : 
                        (N125)? \xz.mem_with_zero_9__20_  : 
                        (N127)? \xz.mem_with_zero_10__20_  : 
                        (N129)? \xz.mem_with_zero_11__20_  : 
                        (N131)? \xz.mem_with_zero_12__20_  : 
                        (N133)? \xz.mem_with_zero_13__20_  : 
                        (N135)? \xz.mem_with_zero_14__20_  : 
                        (N137)? \xz.mem_with_zero_15__20_  : 
                        (N108)? \xz.mem_with_zero_16__20_  : 
                        (N110)? \xz.mem_with_zero_17__20_  : 
                        (N112)? \xz.mem_with_zero_18__20_  : 
                        (N114)? \xz.mem_with_zero_19__20_  : 
                        (N116)? \xz.mem_with_zero_20__20_  : 
                        (N118)? \xz.mem_with_zero_21__20_  : 
                        (N120)? \xz.mem_with_zero_22__20_  : 
                        (N122)? \xz.mem_with_zero_23__20_  : 
                        (N124)? \xz.mem_with_zero_24__20_  : 
                        (N126)? \xz.mem_with_zero_25__20_  : 
                        (N128)? \xz.mem_with_zero_26__20_  : 
                        (N130)? \xz.mem_with_zero_27__20_  : 
                        (N132)? \xz.mem_with_zero_28__20_  : 
                        (N134)? \xz.mem_with_zero_29__20_  : 
                        (N136)? \xz.mem_with_zero_30__20_  : 
                        (N138)? \xz.mem_with_zero_31__20_  : 1'b0;
  assign r_data_o[51] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__19_  : 
                        (N111)? \xz.mem_with_zero_2__19_  : 
                        (N113)? \xz.mem_with_zero_3__19_  : 
                        (N115)? \xz.mem_with_zero_4__19_  : 
                        (N117)? \xz.mem_with_zero_5__19_  : 
                        (N119)? \xz.mem_with_zero_6__19_  : 
                        (N121)? \xz.mem_with_zero_7__19_  : 
                        (N123)? \xz.mem_with_zero_8__19_  : 
                        (N125)? \xz.mem_with_zero_9__19_  : 
                        (N127)? \xz.mem_with_zero_10__19_  : 
                        (N129)? \xz.mem_with_zero_11__19_  : 
                        (N131)? \xz.mem_with_zero_12__19_  : 
                        (N133)? \xz.mem_with_zero_13__19_  : 
                        (N135)? \xz.mem_with_zero_14__19_  : 
                        (N137)? \xz.mem_with_zero_15__19_  : 
                        (N108)? \xz.mem_with_zero_16__19_  : 
                        (N110)? \xz.mem_with_zero_17__19_  : 
                        (N112)? \xz.mem_with_zero_18__19_  : 
                        (N114)? \xz.mem_with_zero_19__19_  : 
                        (N116)? \xz.mem_with_zero_20__19_  : 
                        (N118)? \xz.mem_with_zero_21__19_  : 
                        (N120)? \xz.mem_with_zero_22__19_  : 
                        (N122)? \xz.mem_with_zero_23__19_  : 
                        (N124)? \xz.mem_with_zero_24__19_  : 
                        (N126)? \xz.mem_with_zero_25__19_  : 
                        (N128)? \xz.mem_with_zero_26__19_  : 
                        (N130)? \xz.mem_with_zero_27__19_  : 
                        (N132)? \xz.mem_with_zero_28__19_  : 
                        (N134)? \xz.mem_with_zero_29__19_  : 
                        (N136)? \xz.mem_with_zero_30__19_  : 
                        (N138)? \xz.mem_with_zero_31__19_  : 1'b0;
  assign r_data_o[50] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__18_  : 
                        (N111)? \xz.mem_with_zero_2__18_  : 
                        (N113)? \xz.mem_with_zero_3__18_  : 
                        (N115)? \xz.mem_with_zero_4__18_  : 
                        (N117)? \xz.mem_with_zero_5__18_  : 
                        (N119)? \xz.mem_with_zero_6__18_  : 
                        (N121)? \xz.mem_with_zero_7__18_  : 
                        (N123)? \xz.mem_with_zero_8__18_  : 
                        (N125)? \xz.mem_with_zero_9__18_  : 
                        (N127)? \xz.mem_with_zero_10__18_  : 
                        (N129)? \xz.mem_with_zero_11__18_  : 
                        (N131)? \xz.mem_with_zero_12__18_  : 
                        (N133)? \xz.mem_with_zero_13__18_  : 
                        (N135)? \xz.mem_with_zero_14__18_  : 
                        (N137)? \xz.mem_with_zero_15__18_  : 
                        (N108)? \xz.mem_with_zero_16__18_  : 
                        (N110)? \xz.mem_with_zero_17__18_  : 
                        (N112)? \xz.mem_with_zero_18__18_  : 
                        (N114)? \xz.mem_with_zero_19__18_  : 
                        (N116)? \xz.mem_with_zero_20__18_  : 
                        (N118)? \xz.mem_with_zero_21__18_  : 
                        (N120)? \xz.mem_with_zero_22__18_  : 
                        (N122)? \xz.mem_with_zero_23__18_  : 
                        (N124)? \xz.mem_with_zero_24__18_  : 
                        (N126)? \xz.mem_with_zero_25__18_  : 
                        (N128)? \xz.mem_with_zero_26__18_  : 
                        (N130)? \xz.mem_with_zero_27__18_  : 
                        (N132)? \xz.mem_with_zero_28__18_  : 
                        (N134)? \xz.mem_with_zero_29__18_  : 
                        (N136)? \xz.mem_with_zero_30__18_  : 
                        (N138)? \xz.mem_with_zero_31__18_  : 1'b0;
  assign r_data_o[49] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__17_  : 
                        (N111)? \xz.mem_with_zero_2__17_  : 
                        (N113)? \xz.mem_with_zero_3__17_  : 
                        (N115)? \xz.mem_with_zero_4__17_  : 
                        (N117)? \xz.mem_with_zero_5__17_  : 
                        (N119)? \xz.mem_with_zero_6__17_  : 
                        (N121)? \xz.mem_with_zero_7__17_  : 
                        (N123)? \xz.mem_with_zero_8__17_  : 
                        (N125)? \xz.mem_with_zero_9__17_  : 
                        (N127)? \xz.mem_with_zero_10__17_  : 
                        (N129)? \xz.mem_with_zero_11__17_  : 
                        (N131)? \xz.mem_with_zero_12__17_  : 
                        (N133)? \xz.mem_with_zero_13__17_  : 
                        (N135)? \xz.mem_with_zero_14__17_  : 
                        (N137)? \xz.mem_with_zero_15__17_  : 
                        (N108)? \xz.mem_with_zero_16__17_  : 
                        (N110)? \xz.mem_with_zero_17__17_  : 
                        (N112)? \xz.mem_with_zero_18__17_  : 
                        (N114)? \xz.mem_with_zero_19__17_  : 
                        (N116)? \xz.mem_with_zero_20__17_  : 
                        (N118)? \xz.mem_with_zero_21__17_  : 
                        (N120)? \xz.mem_with_zero_22__17_  : 
                        (N122)? \xz.mem_with_zero_23__17_  : 
                        (N124)? \xz.mem_with_zero_24__17_  : 
                        (N126)? \xz.mem_with_zero_25__17_  : 
                        (N128)? \xz.mem_with_zero_26__17_  : 
                        (N130)? \xz.mem_with_zero_27__17_  : 
                        (N132)? \xz.mem_with_zero_28__17_  : 
                        (N134)? \xz.mem_with_zero_29__17_  : 
                        (N136)? \xz.mem_with_zero_30__17_  : 
                        (N138)? \xz.mem_with_zero_31__17_  : 1'b0;
  assign r_data_o[48] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__16_  : 
                        (N111)? \xz.mem_with_zero_2__16_  : 
                        (N113)? \xz.mem_with_zero_3__16_  : 
                        (N115)? \xz.mem_with_zero_4__16_  : 
                        (N117)? \xz.mem_with_zero_5__16_  : 
                        (N119)? \xz.mem_with_zero_6__16_  : 
                        (N121)? \xz.mem_with_zero_7__16_  : 
                        (N123)? \xz.mem_with_zero_8__16_  : 
                        (N125)? \xz.mem_with_zero_9__16_  : 
                        (N127)? \xz.mem_with_zero_10__16_  : 
                        (N129)? \xz.mem_with_zero_11__16_  : 
                        (N131)? \xz.mem_with_zero_12__16_  : 
                        (N133)? \xz.mem_with_zero_13__16_  : 
                        (N135)? \xz.mem_with_zero_14__16_  : 
                        (N137)? \xz.mem_with_zero_15__16_  : 
                        (N108)? \xz.mem_with_zero_16__16_  : 
                        (N110)? \xz.mem_with_zero_17__16_  : 
                        (N112)? \xz.mem_with_zero_18__16_  : 
                        (N114)? \xz.mem_with_zero_19__16_  : 
                        (N116)? \xz.mem_with_zero_20__16_  : 
                        (N118)? \xz.mem_with_zero_21__16_  : 
                        (N120)? \xz.mem_with_zero_22__16_  : 
                        (N122)? \xz.mem_with_zero_23__16_  : 
                        (N124)? \xz.mem_with_zero_24__16_  : 
                        (N126)? \xz.mem_with_zero_25__16_  : 
                        (N128)? \xz.mem_with_zero_26__16_  : 
                        (N130)? \xz.mem_with_zero_27__16_  : 
                        (N132)? \xz.mem_with_zero_28__16_  : 
                        (N134)? \xz.mem_with_zero_29__16_  : 
                        (N136)? \xz.mem_with_zero_30__16_  : 
                        (N138)? \xz.mem_with_zero_31__16_  : 1'b0;
  assign r_data_o[47] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__15_  : 
                        (N111)? \xz.mem_with_zero_2__15_  : 
                        (N113)? \xz.mem_with_zero_3__15_  : 
                        (N115)? \xz.mem_with_zero_4__15_  : 
                        (N117)? \xz.mem_with_zero_5__15_  : 
                        (N119)? \xz.mem_with_zero_6__15_  : 
                        (N121)? \xz.mem_with_zero_7__15_  : 
                        (N123)? \xz.mem_with_zero_8__15_  : 
                        (N125)? \xz.mem_with_zero_9__15_  : 
                        (N127)? \xz.mem_with_zero_10__15_  : 
                        (N129)? \xz.mem_with_zero_11__15_  : 
                        (N131)? \xz.mem_with_zero_12__15_  : 
                        (N133)? \xz.mem_with_zero_13__15_  : 
                        (N135)? \xz.mem_with_zero_14__15_  : 
                        (N137)? \xz.mem_with_zero_15__15_  : 
                        (N108)? \xz.mem_with_zero_16__15_  : 
                        (N110)? \xz.mem_with_zero_17__15_  : 
                        (N112)? \xz.mem_with_zero_18__15_  : 
                        (N114)? \xz.mem_with_zero_19__15_  : 
                        (N116)? \xz.mem_with_zero_20__15_  : 
                        (N118)? \xz.mem_with_zero_21__15_  : 
                        (N120)? \xz.mem_with_zero_22__15_  : 
                        (N122)? \xz.mem_with_zero_23__15_  : 
                        (N124)? \xz.mem_with_zero_24__15_  : 
                        (N126)? \xz.mem_with_zero_25__15_  : 
                        (N128)? \xz.mem_with_zero_26__15_  : 
                        (N130)? \xz.mem_with_zero_27__15_  : 
                        (N132)? \xz.mem_with_zero_28__15_  : 
                        (N134)? \xz.mem_with_zero_29__15_  : 
                        (N136)? \xz.mem_with_zero_30__15_  : 
                        (N138)? \xz.mem_with_zero_31__15_  : 1'b0;
  assign r_data_o[46] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__14_  : 
                        (N111)? \xz.mem_with_zero_2__14_  : 
                        (N113)? \xz.mem_with_zero_3__14_  : 
                        (N115)? \xz.mem_with_zero_4__14_  : 
                        (N117)? \xz.mem_with_zero_5__14_  : 
                        (N119)? \xz.mem_with_zero_6__14_  : 
                        (N121)? \xz.mem_with_zero_7__14_  : 
                        (N123)? \xz.mem_with_zero_8__14_  : 
                        (N125)? \xz.mem_with_zero_9__14_  : 
                        (N127)? \xz.mem_with_zero_10__14_  : 
                        (N129)? \xz.mem_with_zero_11__14_  : 
                        (N131)? \xz.mem_with_zero_12__14_  : 
                        (N133)? \xz.mem_with_zero_13__14_  : 
                        (N135)? \xz.mem_with_zero_14__14_  : 
                        (N137)? \xz.mem_with_zero_15__14_  : 
                        (N108)? \xz.mem_with_zero_16__14_  : 
                        (N110)? \xz.mem_with_zero_17__14_  : 
                        (N112)? \xz.mem_with_zero_18__14_  : 
                        (N114)? \xz.mem_with_zero_19__14_  : 
                        (N116)? \xz.mem_with_zero_20__14_  : 
                        (N118)? \xz.mem_with_zero_21__14_  : 
                        (N120)? \xz.mem_with_zero_22__14_  : 
                        (N122)? \xz.mem_with_zero_23__14_  : 
                        (N124)? \xz.mem_with_zero_24__14_  : 
                        (N126)? \xz.mem_with_zero_25__14_  : 
                        (N128)? \xz.mem_with_zero_26__14_  : 
                        (N130)? \xz.mem_with_zero_27__14_  : 
                        (N132)? \xz.mem_with_zero_28__14_  : 
                        (N134)? \xz.mem_with_zero_29__14_  : 
                        (N136)? \xz.mem_with_zero_30__14_  : 
                        (N138)? \xz.mem_with_zero_31__14_  : 1'b0;
  assign r_data_o[45] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__13_  : 
                        (N111)? \xz.mem_with_zero_2__13_  : 
                        (N113)? \xz.mem_with_zero_3__13_  : 
                        (N115)? \xz.mem_with_zero_4__13_  : 
                        (N117)? \xz.mem_with_zero_5__13_  : 
                        (N119)? \xz.mem_with_zero_6__13_  : 
                        (N121)? \xz.mem_with_zero_7__13_  : 
                        (N123)? \xz.mem_with_zero_8__13_  : 
                        (N125)? \xz.mem_with_zero_9__13_  : 
                        (N127)? \xz.mem_with_zero_10__13_  : 
                        (N129)? \xz.mem_with_zero_11__13_  : 
                        (N131)? \xz.mem_with_zero_12__13_  : 
                        (N133)? \xz.mem_with_zero_13__13_  : 
                        (N135)? \xz.mem_with_zero_14__13_  : 
                        (N137)? \xz.mem_with_zero_15__13_  : 
                        (N108)? \xz.mem_with_zero_16__13_  : 
                        (N110)? \xz.mem_with_zero_17__13_  : 
                        (N112)? \xz.mem_with_zero_18__13_  : 
                        (N114)? \xz.mem_with_zero_19__13_  : 
                        (N116)? \xz.mem_with_zero_20__13_  : 
                        (N118)? \xz.mem_with_zero_21__13_  : 
                        (N120)? \xz.mem_with_zero_22__13_  : 
                        (N122)? \xz.mem_with_zero_23__13_  : 
                        (N124)? \xz.mem_with_zero_24__13_  : 
                        (N126)? \xz.mem_with_zero_25__13_  : 
                        (N128)? \xz.mem_with_zero_26__13_  : 
                        (N130)? \xz.mem_with_zero_27__13_  : 
                        (N132)? \xz.mem_with_zero_28__13_  : 
                        (N134)? \xz.mem_with_zero_29__13_  : 
                        (N136)? \xz.mem_with_zero_30__13_  : 
                        (N138)? \xz.mem_with_zero_31__13_  : 1'b0;
  assign r_data_o[44] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__12_  : 
                        (N111)? \xz.mem_with_zero_2__12_  : 
                        (N113)? \xz.mem_with_zero_3__12_  : 
                        (N115)? \xz.mem_with_zero_4__12_  : 
                        (N117)? \xz.mem_with_zero_5__12_  : 
                        (N119)? \xz.mem_with_zero_6__12_  : 
                        (N121)? \xz.mem_with_zero_7__12_  : 
                        (N123)? \xz.mem_with_zero_8__12_  : 
                        (N125)? \xz.mem_with_zero_9__12_  : 
                        (N127)? \xz.mem_with_zero_10__12_  : 
                        (N129)? \xz.mem_with_zero_11__12_  : 
                        (N131)? \xz.mem_with_zero_12__12_  : 
                        (N133)? \xz.mem_with_zero_13__12_  : 
                        (N135)? \xz.mem_with_zero_14__12_  : 
                        (N137)? \xz.mem_with_zero_15__12_  : 
                        (N108)? \xz.mem_with_zero_16__12_  : 
                        (N110)? \xz.mem_with_zero_17__12_  : 
                        (N112)? \xz.mem_with_zero_18__12_  : 
                        (N114)? \xz.mem_with_zero_19__12_  : 
                        (N116)? \xz.mem_with_zero_20__12_  : 
                        (N118)? \xz.mem_with_zero_21__12_  : 
                        (N120)? \xz.mem_with_zero_22__12_  : 
                        (N122)? \xz.mem_with_zero_23__12_  : 
                        (N124)? \xz.mem_with_zero_24__12_  : 
                        (N126)? \xz.mem_with_zero_25__12_  : 
                        (N128)? \xz.mem_with_zero_26__12_  : 
                        (N130)? \xz.mem_with_zero_27__12_  : 
                        (N132)? \xz.mem_with_zero_28__12_  : 
                        (N134)? \xz.mem_with_zero_29__12_  : 
                        (N136)? \xz.mem_with_zero_30__12_  : 
                        (N138)? \xz.mem_with_zero_31__12_  : 1'b0;
  assign r_data_o[43] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__11_  : 
                        (N111)? \xz.mem_with_zero_2__11_  : 
                        (N113)? \xz.mem_with_zero_3__11_  : 
                        (N115)? \xz.mem_with_zero_4__11_  : 
                        (N117)? \xz.mem_with_zero_5__11_  : 
                        (N119)? \xz.mem_with_zero_6__11_  : 
                        (N121)? \xz.mem_with_zero_7__11_  : 
                        (N123)? \xz.mem_with_zero_8__11_  : 
                        (N125)? \xz.mem_with_zero_9__11_  : 
                        (N127)? \xz.mem_with_zero_10__11_  : 
                        (N129)? \xz.mem_with_zero_11__11_  : 
                        (N131)? \xz.mem_with_zero_12__11_  : 
                        (N133)? \xz.mem_with_zero_13__11_  : 
                        (N135)? \xz.mem_with_zero_14__11_  : 
                        (N137)? \xz.mem_with_zero_15__11_  : 
                        (N108)? \xz.mem_with_zero_16__11_  : 
                        (N110)? \xz.mem_with_zero_17__11_  : 
                        (N112)? \xz.mem_with_zero_18__11_  : 
                        (N114)? \xz.mem_with_zero_19__11_  : 
                        (N116)? \xz.mem_with_zero_20__11_  : 
                        (N118)? \xz.mem_with_zero_21__11_  : 
                        (N120)? \xz.mem_with_zero_22__11_  : 
                        (N122)? \xz.mem_with_zero_23__11_  : 
                        (N124)? \xz.mem_with_zero_24__11_  : 
                        (N126)? \xz.mem_with_zero_25__11_  : 
                        (N128)? \xz.mem_with_zero_26__11_  : 
                        (N130)? \xz.mem_with_zero_27__11_  : 
                        (N132)? \xz.mem_with_zero_28__11_  : 
                        (N134)? \xz.mem_with_zero_29__11_  : 
                        (N136)? \xz.mem_with_zero_30__11_  : 
                        (N138)? \xz.mem_with_zero_31__11_  : 1'b0;
  assign r_data_o[42] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__10_  : 
                        (N111)? \xz.mem_with_zero_2__10_  : 
                        (N113)? \xz.mem_with_zero_3__10_  : 
                        (N115)? \xz.mem_with_zero_4__10_  : 
                        (N117)? \xz.mem_with_zero_5__10_  : 
                        (N119)? \xz.mem_with_zero_6__10_  : 
                        (N121)? \xz.mem_with_zero_7__10_  : 
                        (N123)? \xz.mem_with_zero_8__10_  : 
                        (N125)? \xz.mem_with_zero_9__10_  : 
                        (N127)? \xz.mem_with_zero_10__10_  : 
                        (N129)? \xz.mem_with_zero_11__10_  : 
                        (N131)? \xz.mem_with_zero_12__10_  : 
                        (N133)? \xz.mem_with_zero_13__10_  : 
                        (N135)? \xz.mem_with_zero_14__10_  : 
                        (N137)? \xz.mem_with_zero_15__10_  : 
                        (N108)? \xz.mem_with_zero_16__10_  : 
                        (N110)? \xz.mem_with_zero_17__10_  : 
                        (N112)? \xz.mem_with_zero_18__10_  : 
                        (N114)? \xz.mem_with_zero_19__10_  : 
                        (N116)? \xz.mem_with_zero_20__10_  : 
                        (N118)? \xz.mem_with_zero_21__10_  : 
                        (N120)? \xz.mem_with_zero_22__10_  : 
                        (N122)? \xz.mem_with_zero_23__10_  : 
                        (N124)? \xz.mem_with_zero_24__10_  : 
                        (N126)? \xz.mem_with_zero_25__10_  : 
                        (N128)? \xz.mem_with_zero_26__10_  : 
                        (N130)? \xz.mem_with_zero_27__10_  : 
                        (N132)? \xz.mem_with_zero_28__10_  : 
                        (N134)? \xz.mem_with_zero_29__10_  : 
                        (N136)? \xz.mem_with_zero_30__10_  : 
                        (N138)? \xz.mem_with_zero_31__10_  : 1'b0;
  assign r_data_o[41] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__9_  : 
                        (N111)? \xz.mem_with_zero_2__9_  : 
                        (N113)? \xz.mem_with_zero_3__9_  : 
                        (N115)? \xz.mem_with_zero_4__9_  : 
                        (N117)? \xz.mem_with_zero_5__9_  : 
                        (N119)? \xz.mem_with_zero_6__9_  : 
                        (N121)? \xz.mem_with_zero_7__9_  : 
                        (N123)? \xz.mem_with_zero_8__9_  : 
                        (N125)? \xz.mem_with_zero_9__9_  : 
                        (N127)? \xz.mem_with_zero_10__9_  : 
                        (N129)? \xz.mem_with_zero_11__9_  : 
                        (N131)? \xz.mem_with_zero_12__9_  : 
                        (N133)? \xz.mem_with_zero_13__9_  : 
                        (N135)? \xz.mem_with_zero_14__9_  : 
                        (N137)? \xz.mem_with_zero_15__9_  : 
                        (N108)? \xz.mem_with_zero_16__9_  : 
                        (N110)? \xz.mem_with_zero_17__9_  : 
                        (N112)? \xz.mem_with_zero_18__9_  : 
                        (N114)? \xz.mem_with_zero_19__9_  : 
                        (N116)? \xz.mem_with_zero_20__9_  : 
                        (N118)? \xz.mem_with_zero_21__9_  : 
                        (N120)? \xz.mem_with_zero_22__9_  : 
                        (N122)? \xz.mem_with_zero_23__9_  : 
                        (N124)? \xz.mem_with_zero_24__9_  : 
                        (N126)? \xz.mem_with_zero_25__9_  : 
                        (N128)? \xz.mem_with_zero_26__9_  : 
                        (N130)? \xz.mem_with_zero_27__9_  : 
                        (N132)? \xz.mem_with_zero_28__9_  : 
                        (N134)? \xz.mem_with_zero_29__9_  : 
                        (N136)? \xz.mem_with_zero_30__9_  : 
                        (N138)? \xz.mem_with_zero_31__9_  : 1'b0;
  assign r_data_o[40] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__8_  : 
                        (N111)? \xz.mem_with_zero_2__8_  : 
                        (N113)? \xz.mem_with_zero_3__8_  : 
                        (N115)? \xz.mem_with_zero_4__8_  : 
                        (N117)? \xz.mem_with_zero_5__8_  : 
                        (N119)? \xz.mem_with_zero_6__8_  : 
                        (N121)? \xz.mem_with_zero_7__8_  : 
                        (N123)? \xz.mem_with_zero_8__8_  : 
                        (N125)? \xz.mem_with_zero_9__8_  : 
                        (N127)? \xz.mem_with_zero_10__8_  : 
                        (N129)? \xz.mem_with_zero_11__8_  : 
                        (N131)? \xz.mem_with_zero_12__8_  : 
                        (N133)? \xz.mem_with_zero_13__8_  : 
                        (N135)? \xz.mem_with_zero_14__8_  : 
                        (N137)? \xz.mem_with_zero_15__8_  : 
                        (N108)? \xz.mem_with_zero_16__8_  : 
                        (N110)? \xz.mem_with_zero_17__8_  : 
                        (N112)? \xz.mem_with_zero_18__8_  : 
                        (N114)? \xz.mem_with_zero_19__8_  : 
                        (N116)? \xz.mem_with_zero_20__8_  : 
                        (N118)? \xz.mem_with_zero_21__8_  : 
                        (N120)? \xz.mem_with_zero_22__8_  : 
                        (N122)? \xz.mem_with_zero_23__8_  : 
                        (N124)? \xz.mem_with_zero_24__8_  : 
                        (N126)? \xz.mem_with_zero_25__8_  : 
                        (N128)? \xz.mem_with_zero_26__8_  : 
                        (N130)? \xz.mem_with_zero_27__8_  : 
                        (N132)? \xz.mem_with_zero_28__8_  : 
                        (N134)? \xz.mem_with_zero_29__8_  : 
                        (N136)? \xz.mem_with_zero_30__8_  : 
                        (N138)? \xz.mem_with_zero_31__8_  : 1'b0;
  assign r_data_o[39] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__7_  : 
                        (N111)? \xz.mem_with_zero_2__7_  : 
                        (N113)? \xz.mem_with_zero_3__7_  : 
                        (N115)? \xz.mem_with_zero_4__7_  : 
                        (N117)? \xz.mem_with_zero_5__7_  : 
                        (N119)? \xz.mem_with_zero_6__7_  : 
                        (N121)? \xz.mem_with_zero_7__7_  : 
                        (N123)? \xz.mem_with_zero_8__7_  : 
                        (N125)? \xz.mem_with_zero_9__7_  : 
                        (N127)? \xz.mem_with_zero_10__7_  : 
                        (N129)? \xz.mem_with_zero_11__7_  : 
                        (N131)? \xz.mem_with_zero_12__7_  : 
                        (N133)? \xz.mem_with_zero_13__7_  : 
                        (N135)? \xz.mem_with_zero_14__7_  : 
                        (N137)? \xz.mem_with_zero_15__7_  : 
                        (N108)? \xz.mem_with_zero_16__7_  : 
                        (N110)? \xz.mem_with_zero_17__7_  : 
                        (N112)? \xz.mem_with_zero_18__7_  : 
                        (N114)? \xz.mem_with_zero_19__7_  : 
                        (N116)? \xz.mem_with_zero_20__7_  : 
                        (N118)? \xz.mem_with_zero_21__7_  : 
                        (N120)? \xz.mem_with_zero_22__7_  : 
                        (N122)? \xz.mem_with_zero_23__7_  : 
                        (N124)? \xz.mem_with_zero_24__7_  : 
                        (N126)? \xz.mem_with_zero_25__7_  : 
                        (N128)? \xz.mem_with_zero_26__7_  : 
                        (N130)? \xz.mem_with_zero_27__7_  : 
                        (N132)? \xz.mem_with_zero_28__7_  : 
                        (N134)? \xz.mem_with_zero_29__7_  : 
                        (N136)? \xz.mem_with_zero_30__7_  : 
                        (N138)? \xz.mem_with_zero_31__7_  : 1'b0;
  assign r_data_o[38] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__6_  : 
                        (N111)? \xz.mem_with_zero_2__6_  : 
                        (N113)? \xz.mem_with_zero_3__6_  : 
                        (N115)? \xz.mem_with_zero_4__6_  : 
                        (N117)? \xz.mem_with_zero_5__6_  : 
                        (N119)? \xz.mem_with_zero_6__6_  : 
                        (N121)? \xz.mem_with_zero_7__6_  : 
                        (N123)? \xz.mem_with_zero_8__6_  : 
                        (N125)? \xz.mem_with_zero_9__6_  : 
                        (N127)? \xz.mem_with_zero_10__6_  : 
                        (N129)? \xz.mem_with_zero_11__6_  : 
                        (N131)? \xz.mem_with_zero_12__6_  : 
                        (N133)? \xz.mem_with_zero_13__6_  : 
                        (N135)? \xz.mem_with_zero_14__6_  : 
                        (N137)? \xz.mem_with_zero_15__6_  : 
                        (N108)? \xz.mem_with_zero_16__6_  : 
                        (N110)? \xz.mem_with_zero_17__6_  : 
                        (N112)? \xz.mem_with_zero_18__6_  : 
                        (N114)? \xz.mem_with_zero_19__6_  : 
                        (N116)? \xz.mem_with_zero_20__6_  : 
                        (N118)? \xz.mem_with_zero_21__6_  : 
                        (N120)? \xz.mem_with_zero_22__6_  : 
                        (N122)? \xz.mem_with_zero_23__6_  : 
                        (N124)? \xz.mem_with_zero_24__6_  : 
                        (N126)? \xz.mem_with_zero_25__6_  : 
                        (N128)? \xz.mem_with_zero_26__6_  : 
                        (N130)? \xz.mem_with_zero_27__6_  : 
                        (N132)? \xz.mem_with_zero_28__6_  : 
                        (N134)? \xz.mem_with_zero_29__6_  : 
                        (N136)? \xz.mem_with_zero_30__6_  : 
                        (N138)? \xz.mem_with_zero_31__6_  : 1'b0;
  assign r_data_o[37] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__5_  : 
                        (N111)? \xz.mem_with_zero_2__5_  : 
                        (N113)? \xz.mem_with_zero_3__5_  : 
                        (N115)? \xz.mem_with_zero_4__5_  : 
                        (N117)? \xz.mem_with_zero_5__5_  : 
                        (N119)? \xz.mem_with_zero_6__5_  : 
                        (N121)? \xz.mem_with_zero_7__5_  : 
                        (N123)? \xz.mem_with_zero_8__5_  : 
                        (N125)? \xz.mem_with_zero_9__5_  : 
                        (N127)? \xz.mem_with_zero_10__5_  : 
                        (N129)? \xz.mem_with_zero_11__5_  : 
                        (N131)? \xz.mem_with_zero_12__5_  : 
                        (N133)? \xz.mem_with_zero_13__5_  : 
                        (N135)? \xz.mem_with_zero_14__5_  : 
                        (N137)? \xz.mem_with_zero_15__5_  : 
                        (N108)? \xz.mem_with_zero_16__5_  : 
                        (N110)? \xz.mem_with_zero_17__5_  : 
                        (N112)? \xz.mem_with_zero_18__5_  : 
                        (N114)? \xz.mem_with_zero_19__5_  : 
                        (N116)? \xz.mem_with_zero_20__5_  : 
                        (N118)? \xz.mem_with_zero_21__5_  : 
                        (N120)? \xz.mem_with_zero_22__5_  : 
                        (N122)? \xz.mem_with_zero_23__5_  : 
                        (N124)? \xz.mem_with_zero_24__5_  : 
                        (N126)? \xz.mem_with_zero_25__5_  : 
                        (N128)? \xz.mem_with_zero_26__5_  : 
                        (N130)? \xz.mem_with_zero_27__5_  : 
                        (N132)? \xz.mem_with_zero_28__5_  : 
                        (N134)? \xz.mem_with_zero_29__5_  : 
                        (N136)? \xz.mem_with_zero_30__5_  : 
                        (N138)? \xz.mem_with_zero_31__5_  : 1'b0;
  assign r_data_o[36] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__4_  : 
                        (N111)? \xz.mem_with_zero_2__4_  : 
                        (N113)? \xz.mem_with_zero_3__4_  : 
                        (N115)? \xz.mem_with_zero_4__4_  : 
                        (N117)? \xz.mem_with_zero_5__4_  : 
                        (N119)? \xz.mem_with_zero_6__4_  : 
                        (N121)? \xz.mem_with_zero_7__4_  : 
                        (N123)? \xz.mem_with_zero_8__4_  : 
                        (N125)? \xz.mem_with_zero_9__4_  : 
                        (N127)? \xz.mem_with_zero_10__4_  : 
                        (N129)? \xz.mem_with_zero_11__4_  : 
                        (N131)? \xz.mem_with_zero_12__4_  : 
                        (N133)? \xz.mem_with_zero_13__4_  : 
                        (N135)? \xz.mem_with_zero_14__4_  : 
                        (N137)? \xz.mem_with_zero_15__4_  : 
                        (N108)? \xz.mem_with_zero_16__4_  : 
                        (N110)? \xz.mem_with_zero_17__4_  : 
                        (N112)? \xz.mem_with_zero_18__4_  : 
                        (N114)? \xz.mem_with_zero_19__4_  : 
                        (N116)? \xz.mem_with_zero_20__4_  : 
                        (N118)? \xz.mem_with_zero_21__4_  : 
                        (N120)? \xz.mem_with_zero_22__4_  : 
                        (N122)? \xz.mem_with_zero_23__4_  : 
                        (N124)? \xz.mem_with_zero_24__4_  : 
                        (N126)? \xz.mem_with_zero_25__4_  : 
                        (N128)? \xz.mem_with_zero_26__4_  : 
                        (N130)? \xz.mem_with_zero_27__4_  : 
                        (N132)? \xz.mem_with_zero_28__4_  : 
                        (N134)? \xz.mem_with_zero_29__4_  : 
                        (N136)? \xz.mem_with_zero_30__4_  : 
                        (N138)? \xz.mem_with_zero_31__4_  : 1'b0;
  assign r_data_o[35] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__3_  : 
                        (N111)? \xz.mem_with_zero_2__3_  : 
                        (N113)? \xz.mem_with_zero_3__3_  : 
                        (N115)? \xz.mem_with_zero_4__3_  : 
                        (N117)? \xz.mem_with_zero_5__3_  : 
                        (N119)? \xz.mem_with_zero_6__3_  : 
                        (N121)? \xz.mem_with_zero_7__3_  : 
                        (N123)? \xz.mem_with_zero_8__3_  : 
                        (N125)? \xz.mem_with_zero_9__3_  : 
                        (N127)? \xz.mem_with_zero_10__3_  : 
                        (N129)? \xz.mem_with_zero_11__3_  : 
                        (N131)? \xz.mem_with_zero_12__3_  : 
                        (N133)? \xz.mem_with_zero_13__3_  : 
                        (N135)? \xz.mem_with_zero_14__3_  : 
                        (N137)? \xz.mem_with_zero_15__3_  : 
                        (N108)? \xz.mem_with_zero_16__3_  : 
                        (N110)? \xz.mem_with_zero_17__3_  : 
                        (N112)? \xz.mem_with_zero_18__3_  : 
                        (N114)? \xz.mem_with_zero_19__3_  : 
                        (N116)? \xz.mem_with_zero_20__3_  : 
                        (N118)? \xz.mem_with_zero_21__3_  : 
                        (N120)? \xz.mem_with_zero_22__3_  : 
                        (N122)? \xz.mem_with_zero_23__3_  : 
                        (N124)? \xz.mem_with_zero_24__3_  : 
                        (N126)? \xz.mem_with_zero_25__3_  : 
                        (N128)? \xz.mem_with_zero_26__3_  : 
                        (N130)? \xz.mem_with_zero_27__3_  : 
                        (N132)? \xz.mem_with_zero_28__3_  : 
                        (N134)? \xz.mem_with_zero_29__3_  : 
                        (N136)? \xz.mem_with_zero_30__3_  : 
                        (N138)? \xz.mem_with_zero_31__3_  : 1'b0;
  assign r_data_o[34] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__2_  : 
                        (N111)? \xz.mem_with_zero_2__2_  : 
                        (N113)? \xz.mem_with_zero_3__2_  : 
                        (N115)? \xz.mem_with_zero_4__2_  : 
                        (N117)? \xz.mem_with_zero_5__2_  : 
                        (N119)? \xz.mem_with_zero_6__2_  : 
                        (N121)? \xz.mem_with_zero_7__2_  : 
                        (N123)? \xz.mem_with_zero_8__2_  : 
                        (N125)? \xz.mem_with_zero_9__2_  : 
                        (N127)? \xz.mem_with_zero_10__2_  : 
                        (N129)? \xz.mem_with_zero_11__2_  : 
                        (N131)? \xz.mem_with_zero_12__2_  : 
                        (N133)? \xz.mem_with_zero_13__2_  : 
                        (N135)? \xz.mem_with_zero_14__2_  : 
                        (N137)? \xz.mem_with_zero_15__2_  : 
                        (N108)? \xz.mem_with_zero_16__2_  : 
                        (N110)? \xz.mem_with_zero_17__2_  : 
                        (N112)? \xz.mem_with_zero_18__2_  : 
                        (N114)? \xz.mem_with_zero_19__2_  : 
                        (N116)? \xz.mem_with_zero_20__2_  : 
                        (N118)? \xz.mem_with_zero_21__2_  : 
                        (N120)? \xz.mem_with_zero_22__2_  : 
                        (N122)? \xz.mem_with_zero_23__2_  : 
                        (N124)? \xz.mem_with_zero_24__2_  : 
                        (N126)? \xz.mem_with_zero_25__2_  : 
                        (N128)? \xz.mem_with_zero_26__2_  : 
                        (N130)? \xz.mem_with_zero_27__2_  : 
                        (N132)? \xz.mem_with_zero_28__2_  : 
                        (N134)? \xz.mem_with_zero_29__2_  : 
                        (N136)? \xz.mem_with_zero_30__2_  : 
                        (N138)? \xz.mem_with_zero_31__2_  : 1'b0;
  assign r_data_o[33] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__1_  : 
                        (N111)? \xz.mem_with_zero_2__1_  : 
                        (N113)? \xz.mem_with_zero_3__1_  : 
                        (N115)? \xz.mem_with_zero_4__1_  : 
                        (N117)? \xz.mem_with_zero_5__1_  : 
                        (N119)? \xz.mem_with_zero_6__1_  : 
                        (N121)? \xz.mem_with_zero_7__1_  : 
                        (N123)? \xz.mem_with_zero_8__1_  : 
                        (N125)? \xz.mem_with_zero_9__1_  : 
                        (N127)? \xz.mem_with_zero_10__1_  : 
                        (N129)? \xz.mem_with_zero_11__1_  : 
                        (N131)? \xz.mem_with_zero_12__1_  : 
                        (N133)? \xz.mem_with_zero_13__1_  : 
                        (N135)? \xz.mem_with_zero_14__1_  : 
                        (N137)? \xz.mem_with_zero_15__1_  : 
                        (N108)? \xz.mem_with_zero_16__1_  : 
                        (N110)? \xz.mem_with_zero_17__1_  : 
                        (N112)? \xz.mem_with_zero_18__1_  : 
                        (N114)? \xz.mem_with_zero_19__1_  : 
                        (N116)? \xz.mem_with_zero_20__1_  : 
                        (N118)? \xz.mem_with_zero_21__1_  : 
                        (N120)? \xz.mem_with_zero_22__1_  : 
                        (N122)? \xz.mem_with_zero_23__1_  : 
                        (N124)? \xz.mem_with_zero_24__1_  : 
                        (N126)? \xz.mem_with_zero_25__1_  : 
                        (N128)? \xz.mem_with_zero_26__1_  : 
                        (N130)? \xz.mem_with_zero_27__1_  : 
                        (N132)? \xz.mem_with_zero_28__1_  : 
                        (N134)? \xz.mem_with_zero_29__1_  : 
                        (N136)? \xz.mem_with_zero_30__1_  : 
                        (N138)? \xz.mem_with_zero_31__1_  : 1'b0;
  assign r_data_o[32] = (N107)? 1'b0 : 
                        (N109)? \xz.mem_with_zero_1__0_  : 
                        (N111)? \xz.mem_with_zero_2__0_  : 
                        (N113)? \xz.mem_with_zero_3__0_  : 
                        (N115)? \xz.mem_with_zero_4__0_  : 
                        (N117)? \xz.mem_with_zero_5__0_  : 
                        (N119)? \xz.mem_with_zero_6__0_  : 
                        (N121)? \xz.mem_with_zero_7__0_  : 
                        (N123)? \xz.mem_with_zero_8__0_  : 
                        (N125)? \xz.mem_with_zero_9__0_  : 
                        (N127)? \xz.mem_with_zero_10__0_  : 
                        (N129)? \xz.mem_with_zero_11__0_  : 
                        (N131)? \xz.mem_with_zero_12__0_  : 
                        (N133)? \xz.mem_with_zero_13__0_  : 
                        (N135)? \xz.mem_with_zero_14__0_  : 
                        (N137)? \xz.mem_with_zero_15__0_  : 
                        (N108)? \xz.mem_with_zero_16__0_  : 
                        (N110)? \xz.mem_with_zero_17__0_  : 
                        (N112)? \xz.mem_with_zero_18__0_  : 
                        (N114)? \xz.mem_with_zero_19__0_  : 
                        (N116)? \xz.mem_with_zero_20__0_  : 
                        (N118)? \xz.mem_with_zero_21__0_  : 
                        (N120)? \xz.mem_with_zero_22__0_  : 
                        (N122)? \xz.mem_with_zero_23__0_  : 
                        (N124)? \xz.mem_with_zero_24__0_  : 
                        (N126)? \xz.mem_with_zero_25__0_  : 
                        (N128)? \xz.mem_with_zero_26__0_  : 
                        (N130)? \xz.mem_with_zero_27__0_  : 
                        (N132)? \xz.mem_with_zero_28__0_  : 
                        (N134)? \xz.mem_with_zero_29__0_  : 
                        (N136)? \xz.mem_with_zero_30__0_  : 
                        (N138)? \xz.mem_with_zero_31__0_  : 1'b0;
  assign N203 = w_addr_i[3] | w_addr_i[4];
  assign N204 = w_addr_i[2] | N203;
  assign N205 = w_addr_i[1] | N204;
  assign N206 = w_addr_i[0] | N205;
  assign N207 = w_addr_i[3] & w_addr_i[4];
  assign N208 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N209 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N210 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N211 = ~w_addr_i[2];
  assign N212 = w_addr_i[0] & w_addr_i[1];
  assign N213 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N214 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N215 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N216 = w_addr_i[2] & N212;
  assign N217 = w_addr_i[2] & N213;
  assign N218 = w_addr_i[2] & N214;
  assign N219 = w_addr_i[2] & N215;
  assign N220 = N211 & N212;
  assign N221 = N211 & N213;
  assign N222 = N211 & N214;
  assign N223 = N211 & N215;
  assign N171 = N207 & N216;
  assign N170 = N207 & N217;
  assign N169 = N207 & N218;
  assign N168 = N207 & N219;
  assign N167 = N207 & N220;
  assign N166 = N207 & N221;
  assign N165 = N207 & N222;
  assign N164 = N207 & N223;
  assign N163 = N208 & N216;
  assign N162 = N208 & N217;
  assign N161 = N208 & N218;
  assign N160 = N208 & N219;
  assign N159 = N208 & N220;
  assign N158 = N208 & N221;
  assign N157 = N208 & N222;
  assign N156 = N208 & N223;
  assign N155 = N209 & N216;
  assign N154 = N209 & N217;
  assign N153 = N209 & N218;
  assign N152 = N209 & N219;
  assign N151 = N209 & N220;
  assign N150 = N209 & N221;
  assign N149 = N209 & N222;
  assign N148 = N209 & N223;
  assign N147 = N210 & N216;
  assign N146 = N210 & N217;
  assign N145 = N210 & N218;
  assign N144 = N210 & N219;
  assign N143 = N210 & N220;
  assign N142 = N210 & N221;
  assign N141 = N210 & N222;
  assign { N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172 } = (N8)? { N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } : 
                                                                                                                                                                                                        (N140)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N139;
  assign N9 = ~r_addr_r[0];
  assign N10 = ~r_addr_r[1];
  assign N11 = N9 & N10;
  assign N12 = N9 & r_addr_r[1];
  assign N13 = r_addr_r[0] & N10;
  assign N14 = r_addr_r[0] & r_addr_r[1];
  assign N15 = ~r_addr_r[2];
  assign N16 = N11 & N15;
  assign N17 = N11 & r_addr_r[2];
  assign N18 = N13 & N15;
  assign N19 = N13 & r_addr_r[2];
  assign N20 = N12 & N15;
  assign N21 = N12 & r_addr_r[2];
  assign N22 = N14 & N15;
  assign N23 = N14 & r_addr_r[2];
  assign N24 = ~r_addr_r[3];
  assign N25 = N16 & N24;
  assign N26 = N16 & r_addr_r[3];
  assign N27 = N18 & N24;
  assign N28 = N18 & r_addr_r[3];
  assign N29 = N20 & N24;
  assign N30 = N20 & r_addr_r[3];
  assign N31 = N22 & N24;
  assign N32 = N22 & r_addr_r[3];
  assign N33 = N17 & N24;
  assign N34 = N17 & r_addr_r[3];
  assign N35 = N19 & N24;
  assign N36 = N19 & r_addr_r[3];
  assign N37 = N21 & N24;
  assign N38 = N21 & r_addr_r[3];
  assign N39 = N23 & N24;
  assign N40 = N23 & r_addr_r[3];
  assign N41 = ~r_addr_r[4];
  assign N42 = N25 & N41;
  assign N43 = N25 & r_addr_r[4];
  assign N44 = N27 & N41;
  assign N45 = N27 & r_addr_r[4];
  assign N46 = N29 & N41;
  assign N47 = N29 & r_addr_r[4];
  assign N48 = N31 & N41;
  assign N49 = N31 & r_addr_r[4];
  assign N50 = N33 & N41;
  assign N51 = N33 & r_addr_r[4];
  assign N52 = N35 & N41;
  assign N53 = N35 & r_addr_r[4];
  assign N54 = N37 & N41;
  assign N55 = N37 & r_addr_r[4];
  assign N56 = N39 & N41;
  assign N57 = N39 & r_addr_r[4];
  assign N58 = N26 & N41;
  assign N59 = N26 & r_addr_r[4];
  assign N60 = N28 & N41;
  assign N61 = N28 & r_addr_r[4];
  assign N62 = N30 & N41;
  assign N63 = N30 & r_addr_r[4];
  assign N64 = N32 & N41;
  assign N65 = N32 & r_addr_r[4];
  assign N66 = N34 & N41;
  assign N67 = N34 & r_addr_r[4];
  assign N68 = N36 & N41;
  assign N69 = N36 & r_addr_r[4];
  assign N70 = N38 & N41;
  assign N71 = N38 & r_addr_r[4];
  assign N72 = N40 & N41;
  assign N73 = N40 & r_addr_r[4];
  assign N74 = ~r_addr_r[5];
  assign N75 = ~r_addr_r[6];
  assign N76 = N74 & N75;
  assign N77 = N74 & r_addr_r[6];
  assign N78 = r_addr_r[5] & N75;
  assign N79 = r_addr_r[5] & r_addr_r[6];
  assign N80 = ~r_addr_r[7];
  assign N81 = N76 & N80;
  assign N82 = N76 & r_addr_r[7];
  assign N83 = N78 & N80;
  assign N84 = N78 & r_addr_r[7];
  assign N85 = N77 & N80;
  assign N86 = N77 & r_addr_r[7];
  assign N87 = N79 & N80;
  assign N88 = N79 & r_addr_r[7];
  assign N89 = ~r_addr_r[8];
  assign N90 = N81 & N89;
  assign N91 = N81 & r_addr_r[8];
  assign N92 = N83 & N89;
  assign N93 = N83 & r_addr_r[8];
  assign N94 = N85 & N89;
  assign N95 = N85 & r_addr_r[8];
  assign N96 = N87 & N89;
  assign N97 = N87 & r_addr_r[8];
  assign N98 = N82 & N89;
  assign N99 = N82 & r_addr_r[8];
  assign N100 = N84 & N89;
  assign N101 = N84 & r_addr_r[8];
  assign N102 = N86 & N89;
  assign N103 = N86 & r_addr_r[8];
  assign N104 = N88 & N89;
  assign N105 = N88 & r_addr_r[8];
  assign N106 = ~r_addr_r[9];
  assign N107 = N90 & N106;
  assign N108 = N90 & r_addr_r[9];
  assign N109 = N92 & N106;
  assign N110 = N92 & r_addr_r[9];
  assign N111 = N94 & N106;
  assign N112 = N94 & r_addr_r[9];
  assign N113 = N96 & N106;
  assign N114 = N96 & r_addr_r[9];
  assign N115 = N98 & N106;
  assign N116 = N98 & r_addr_r[9];
  assign N117 = N100 & N106;
  assign N118 = N100 & r_addr_r[9];
  assign N119 = N102 & N106;
  assign N120 = N102 & r_addr_r[9];
  assign N121 = N104 & N106;
  assign N122 = N104 & r_addr_r[9];
  assign N123 = N91 & N106;
  assign N124 = N91 & r_addr_r[9];
  assign N125 = N93 & N106;
  assign N126 = N93 & r_addr_r[9];
  assign N127 = N95 & N106;
  assign N128 = N95 & r_addr_r[9];
  assign N129 = N97 & N106;
  assign N130 = N97 & r_addr_r[9];
  assign N131 = N99 & N106;
  assign N132 = N99 & r_addr_r[9];
  assign N133 = N101 & N106;
  assign N134 = N101 & r_addr_r[9];
  assign N135 = N103 & N106;
  assign N136 = N103 & r_addr_r[9];
  assign N137 = N105 & N106;
  assign N138 = N105 & r_addr_r[9];
  assign N139 = w_v_i & N206;
  assign N140 = ~N139;

  always @(posedge clk_i) begin
    if(r_v_i[1]) begin
      r_addr_r_9_sv2v_reg <= r_addr_i[9];
      r_addr_r_8_sv2v_reg <= r_addr_i[8];
      r_addr_r_7_sv2v_reg <= r_addr_i[7];
      r_addr_r_6_sv2v_reg <= r_addr_i[6];
      r_addr_r_5_sv2v_reg <= r_addr_i[5];
    end 
    if(r_v_i[0]) begin
      r_addr_r_4_sv2v_reg <= r_addr_i[4];
      r_addr_r_3_sv2v_reg <= r_addr_i[3];
      r_addr_r_2_sv2v_reg <= r_addr_i[2];
      r_addr_r_1_sv2v_reg <= r_addr_i[1];
      r_addr_r_0_sv2v_reg <= r_addr_i[0];
    end 
    if(N202) begin
      \xz.mem_with_zero_31__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_31__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_31__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_31__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_31__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_31__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_31__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_31__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_31__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_31__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_31__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_31__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_31__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_31__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_31__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_31__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_31__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_31__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_31__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_31__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_31__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_31__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_31__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_31__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_31__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_31__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_31__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_31__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_31__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_31__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_31__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_31__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N201) begin
      \xz.mem_with_zero_30__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_30__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_30__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_30__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_30__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_30__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_30__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_30__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_30__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_30__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_30__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_30__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_30__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_30__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_30__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_30__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_30__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_30__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_30__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_30__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_30__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_30__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_30__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_30__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_30__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_30__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_30__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_30__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_30__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_30__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_30__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_30__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N200) begin
      \xz.mem_with_zero_29__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_29__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_29__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_29__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_29__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_29__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_29__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_29__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_29__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_29__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_29__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_29__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_29__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_29__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_29__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_29__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_29__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_29__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_29__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_29__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_29__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_29__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_29__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_29__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_29__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_29__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_29__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_29__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_29__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_29__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_29__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_29__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N199) begin
      \xz.mem_with_zero_28__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_28__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_28__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_28__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_28__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_28__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_28__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_28__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_28__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_28__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_28__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_28__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_28__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_28__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_28__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_28__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_28__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_28__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_28__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_28__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_28__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_28__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_28__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_28__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_28__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_28__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_28__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_28__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_28__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_28__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_28__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_28__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N198) begin
      \xz.mem_with_zero_27__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_27__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_27__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_27__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_27__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_27__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_27__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_27__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_27__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_27__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_27__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_27__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_27__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_27__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_27__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_27__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_27__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_27__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_27__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_27__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_27__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_27__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_27__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_27__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_27__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_27__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_27__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_27__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_27__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_27__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_27__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_27__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N197) begin
      \xz.mem_with_zero_26__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_26__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_26__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_26__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_26__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_26__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_26__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_26__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_26__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_26__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_26__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_26__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_26__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_26__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_26__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_26__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_26__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_26__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_26__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_26__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_26__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_26__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_26__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_26__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_26__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_26__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_26__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_26__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_26__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_26__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_26__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_26__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N196) begin
      \xz.mem_with_zero_25__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_25__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_25__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_25__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_25__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_25__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_25__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_25__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_25__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_25__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_25__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_25__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_25__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_25__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_25__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_25__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_25__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_25__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_25__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_25__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_25__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_25__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_25__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_25__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_25__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_25__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_25__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_25__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_25__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_25__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_25__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_25__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N195) begin
      \xz.mem_with_zero_24__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_24__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_24__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_24__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_24__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_24__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_24__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_24__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_24__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_24__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_24__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_24__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_24__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_24__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_24__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_24__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_24__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_24__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_24__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_24__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_24__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_24__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_24__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_24__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_24__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_24__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_24__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_24__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_24__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_24__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_24__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_24__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N194) begin
      \xz.mem_with_zero_23__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_23__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_23__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_23__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_23__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_23__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_23__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_23__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_23__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_23__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_23__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_23__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_23__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_23__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_23__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_23__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_23__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_23__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_23__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_23__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_23__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_23__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_23__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_23__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_23__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_23__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_23__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_23__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_23__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_23__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_23__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_23__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N193) begin
      \xz.mem_with_zero_22__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_22__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_22__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_22__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_22__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_22__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_22__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_22__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_22__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_22__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_22__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_22__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_22__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_22__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_22__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_22__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_22__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_22__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_22__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_22__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_22__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_22__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_22__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_22__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_22__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_22__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_22__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_22__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_22__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_22__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_22__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_22__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N192) begin
      \xz.mem_with_zero_21__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_21__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_21__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_21__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_21__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_21__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_21__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_21__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_21__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_21__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_21__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_21__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_21__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_21__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_21__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_21__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_21__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_21__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_21__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_21__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_21__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_21__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_21__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_21__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_21__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_21__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_21__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_21__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_21__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_21__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_21__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_21__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N191) begin
      \xz.mem_with_zero_20__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_20__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_20__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_20__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_20__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_20__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_20__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_20__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_20__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_20__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_20__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_20__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_20__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_20__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_20__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_20__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_20__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_20__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_20__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_20__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_20__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_20__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_20__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_20__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_20__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_20__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_20__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_20__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_20__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_20__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_20__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_20__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N190) begin
      \xz.mem_with_zero_19__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_19__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_19__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_19__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_19__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_19__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_19__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_19__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_19__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_19__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_19__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_19__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_19__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_19__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_19__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_19__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_19__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_19__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_19__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_19__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_19__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_19__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_19__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_19__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_19__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_19__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_19__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_19__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_19__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_19__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_19__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_19__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N189) begin
      \xz.mem_with_zero_18__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_18__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_18__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_18__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_18__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_18__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_18__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_18__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_18__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_18__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_18__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_18__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_18__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_18__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_18__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_18__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_18__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_18__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_18__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_18__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_18__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_18__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_18__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_18__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_18__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_18__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_18__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_18__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_18__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_18__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_18__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_18__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N188) begin
      \xz.mem_with_zero_17__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_17__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_17__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_17__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_17__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_17__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_17__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_17__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_17__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_17__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_17__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_17__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_17__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_17__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_17__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_17__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_17__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_17__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_17__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_17__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_17__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_17__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_17__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_17__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_17__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_17__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_17__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_17__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_17__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_17__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_17__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_17__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N187) begin
      \xz.mem_with_zero_16__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_16__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_16__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_16__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_16__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_16__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_16__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_16__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_16__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_16__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_16__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_16__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_16__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_16__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_16__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_16__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_16__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_16__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_16__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_16__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_16__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_16__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_16__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_16__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_16__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_16__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_16__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_16__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_16__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_16__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_16__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_16__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N186) begin
      \xz.mem_with_zero_15__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_15__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_15__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_15__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_15__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_15__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_15__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_15__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_15__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_15__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_15__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_15__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_15__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_15__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_15__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_15__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_15__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_15__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_15__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_15__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_15__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_15__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_15__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_15__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_15__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_15__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_15__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_15__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_15__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_15__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_15__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_15__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N185) begin
      \xz.mem_with_zero_14__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_14__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_14__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_14__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_14__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_14__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_14__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_14__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_14__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_14__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_14__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_14__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_14__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_14__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_14__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_14__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_14__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_14__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_14__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_14__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_14__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_14__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_14__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_14__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_14__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_14__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_14__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_14__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_14__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_14__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_14__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_14__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N184) begin
      \xz.mem_with_zero_13__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_13__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_13__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_13__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_13__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_13__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_13__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_13__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_13__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_13__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_13__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_13__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_13__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_13__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_13__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_13__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_13__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_13__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_13__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_13__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_13__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_13__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_13__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_13__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_13__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_13__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_13__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_13__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_13__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_13__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_13__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_13__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N183) begin
      \xz.mem_with_zero_12__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_12__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_12__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_12__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_12__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_12__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_12__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_12__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_12__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_12__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_12__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_12__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_12__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_12__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_12__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_12__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_12__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_12__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_12__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_12__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_12__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_12__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_12__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_12__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_12__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_12__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_12__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_12__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_12__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_12__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_12__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_12__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N182) begin
      \xz.mem_with_zero_11__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_11__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_11__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_11__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_11__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_11__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_11__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_11__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_11__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_11__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_11__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_11__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_11__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_11__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_11__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_11__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_11__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_11__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_11__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_11__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_11__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_11__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_11__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_11__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_11__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_11__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_11__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_11__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_11__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_11__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_11__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_11__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N181) begin
      \xz.mem_with_zero_10__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_10__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_10__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_10__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_10__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_10__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_10__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_10__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_10__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_10__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_10__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_10__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_10__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_10__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_10__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_10__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_10__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_10__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_10__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_10__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_10__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_10__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_10__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_10__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_10__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_10__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_10__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_10__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_10__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_10__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_10__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_10__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N180) begin
      \xz.mem_with_zero_9__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_9__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_9__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_9__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_9__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_9__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_9__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_9__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_9__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_9__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_9__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_9__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_9__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_9__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_9__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_9__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_9__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_9__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_9__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_9__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_9__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_9__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_9__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_9__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_9__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_9__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_9__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_9__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_9__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_9__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_9__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_9__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N179) begin
      \xz.mem_with_zero_8__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_8__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_8__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_8__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_8__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_8__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_8__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_8__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_8__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_8__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_8__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_8__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_8__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_8__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_8__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_8__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_8__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_8__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_8__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_8__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_8__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_8__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_8__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_8__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_8__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_8__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_8__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_8__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_8__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_8__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_8__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_8__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N178) begin
      \xz.mem_with_zero_7__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_7__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_7__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_7__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_7__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_7__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_7__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_7__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_7__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_7__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_7__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_7__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_7__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_7__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_7__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_7__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_7__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_7__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_7__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_7__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_7__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_7__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_7__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_7__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_7__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_7__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_7__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_7__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_7__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_7__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_7__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_7__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N177) begin
      \xz.mem_with_zero_6__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_6__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_6__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_6__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_6__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_6__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_6__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_6__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_6__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_6__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_6__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_6__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_6__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_6__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_6__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_6__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_6__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_6__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_6__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_6__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_6__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_6__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_6__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_6__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_6__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_6__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_6__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_6__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_6__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_6__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_6__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_6__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N176) begin
      \xz.mem_with_zero_5__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_5__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_5__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_5__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_5__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_5__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_5__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_5__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_5__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_5__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_5__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_5__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_5__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_5__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_5__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_5__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_5__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_5__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_5__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_5__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_5__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_5__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_5__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_5__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_5__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_5__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_5__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_5__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_5__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_5__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_5__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_5__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N175) begin
      \xz.mem_with_zero_4__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_4__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_4__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_4__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_4__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_4__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_4__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_4__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_4__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_4__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_4__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_4__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_4__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_4__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_4__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_4__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_4__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_4__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_4__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_4__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_4__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_4__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_4__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_4__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_4__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_4__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_4__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_4__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_4__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_4__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_4__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_4__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N174) begin
      \xz.mem_with_zero_3__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_3__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_3__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_3__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_3__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_3__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_3__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_3__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_3__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_3__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_3__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_3__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_3__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_3__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_3__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_3__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_3__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_3__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_3__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_3__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_3__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_3__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_3__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_3__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_3__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_3__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_3__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_3__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_3__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_3__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_3__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_3__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N173) begin
      \xz.mem_with_zero_2__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_2__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_2__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_2__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_2__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_2__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_2__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_2__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_2__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_2__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_2__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_2__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_2__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_2__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_2__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_2__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_2__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_2__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_2__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_2__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_2__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_2__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_2__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_2__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_2__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_2__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_2__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_2__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_2__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_2__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_2__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_2__0__sv2v_reg  <= w_data_i[0];
    end 
    if(N172) begin
      \xz.mem_with_zero_1__31__sv2v_reg  <= w_data_i[31];
      \xz.mem_with_zero_1__30__sv2v_reg  <= w_data_i[30];
      \xz.mem_with_zero_1__29__sv2v_reg  <= w_data_i[29];
      \xz.mem_with_zero_1__28__sv2v_reg  <= w_data_i[28];
      \xz.mem_with_zero_1__27__sv2v_reg  <= w_data_i[27];
      \xz.mem_with_zero_1__26__sv2v_reg  <= w_data_i[26];
      \xz.mem_with_zero_1__25__sv2v_reg  <= w_data_i[25];
      \xz.mem_with_zero_1__24__sv2v_reg  <= w_data_i[24];
      \xz.mem_with_zero_1__23__sv2v_reg  <= w_data_i[23];
      \xz.mem_with_zero_1__22__sv2v_reg  <= w_data_i[22];
      \xz.mem_with_zero_1__21__sv2v_reg  <= w_data_i[21];
      \xz.mem_with_zero_1__20__sv2v_reg  <= w_data_i[20];
      \xz.mem_with_zero_1__19__sv2v_reg  <= w_data_i[19];
      \xz.mem_with_zero_1__18__sv2v_reg  <= w_data_i[18];
      \xz.mem_with_zero_1__17__sv2v_reg  <= w_data_i[17];
      \xz.mem_with_zero_1__16__sv2v_reg  <= w_data_i[16];
      \xz.mem_with_zero_1__15__sv2v_reg  <= w_data_i[15];
      \xz.mem_with_zero_1__14__sv2v_reg  <= w_data_i[14];
      \xz.mem_with_zero_1__13__sv2v_reg  <= w_data_i[13];
      \xz.mem_with_zero_1__12__sv2v_reg  <= w_data_i[12];
      \xz.mem_with_zero_1__11__sv2v_reg  <= w_data_i[11];
      \xz.mem_with_zero_1__10__sv2v_reg  <= w_data_i[10];
      \xz.mem_with_zero_1__9__sv2v_reg  <= w_data_i[9];
      \xz.mem_with_zero_1__8__sv2v_reg  <= w_data_i[8];
      \xz.mem_with_zero_1__7__sv2v_reg  <= w_data_i[7];
      \xz.mem_with_zero_1__6__sv2v_reg  <= w_data_i[6];
      \xz.mem_with_zero_1__5__sv2v_reg  <= w_data_i[5];
      \xz.mem_with_zero_1__4__sv2v_reg  <= w_data_i[4];
      \xz.mem_with_zero_1__3__sv2v_reg  <= w_data_i[3];
      \xz.mem_with_zero_1__2__sv2v_reg  <= w_data_i[2];
      \xz.mem_with_zero_1__1__sv2v_reg  <= w_data_i[1];
      \xz.mem_with_zero_1__0__sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module regfile_width_p32_els_p32_num_rs_p2_x0_tied_to_zero_p1
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [4:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_v_i;
  input [9:0] r_addr_i;
  output [63:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  wire [63:0] r_data_o;

  regfile_synth_width_p32_els_p32_num_rs_p2_x0_tied_to_zero_p1
  \synth.rf 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_transpose_width_p32_els_p1
(
  i,
  o
);

  input [31:0] i;
  output [31:0] o;
  wire [31:0] o;
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_decode_num_out_p32
(
  i,
  o
);

  input [4:0] i;
  output [31:0] o;
  wire [31:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_decode_with_v_num_out_p32
(
  i,
  v_i,
  o
);

  input [4:0] i;
  output [31:0] o;
  input v_i;
  wire [31:0] o,lo;

  bsg_decode_num_out_p32
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[31] = v_i & lo[31];
  assign o[30] = v_i & lo[30];
  assign o[29] = v_i & lo[29];
  assign o[28] = v_i & lo[28];
  assign o[27] = v_i & lo[27];
  assign o[26] = v_i & lo[26];
  assign o[25] = v_i & lo[25];
  assign o[24] = v_i & lo[24];
  assign o[23] = v_i & lo[23];
  assign o[22] = v_i & lo[22];
  assign o[21] = v_i & lo[21];
  assign o[20] = v_i & lo[20];
  assign o[19] = v_i & lo[19];
  assign o[18] = v_i & lo[18];
  assign o[17] = v_i & lo[17];
  assign o[16] = v_i & lo[16];
  assign o[15] = v_i & lo[15];
  assign o[14] = v_i & lo[14];
  assign o[13] = v_i & lo[13];
  assign o[12] = v_i & lo[12];
  assign o[11] = v_i & lo[11];
  assign o[10] = v_i & lo[10];
  assign o[9] = v_i & lo[9];
  assign o[8] = v_i & lo[8];
  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_transpose_width_p2_els_p1
(
  i,
  o
);

  input [1:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module scoreboard_els_p32_num_src_port_p2_num_clear_port_p1_x0_tied_to_zero_p1
(
  clk_i,
  reset_i,
  src_id_i,
  dest_id_i,
  op_reads_rf_i,
  op_writes_rf_i,
  score_i,
  score_id_i,
  clear_i,
  clear_id_i,
  dependency_o
);

  input [9:0] src_id_i;
  input [4:0] dest_id_i;
  input [1:0] op_reads_rf_i;
  input [4:0] score_id_i;
  input [0:0] clear_i;
  input [4:0] clear_id_i;
  input clk_i;
  input reset_i;
  input op_writes_rf_i;
  input score_i;
  output dependency_o;
  wire dependency_o,_0_net_,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,rd_depend_on_sb,N198,N199,N200,N201,N202,N203,
  rd_depend_on_score,depend_on_sb,depend_on_score,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217;
  wire [31:0] clear_by_port,clear_by_port_t,score_bits,scoreboard_r;
  wire [1:0] rs_depend_on_sb,rs_on_clear,rs_on_clear_t,rs_depend_on_score;
  wire [0:0] rd_on_clear;
  reg scoreboard_r_31_sv2v_reg,scoreboard_r_30_sv2v_reg,scoreboard_r_29_sv2v_reg,
  scoreboard_r_28_sv2v_reg,scoreboard_r_27_sv2v_reg,scoreboard_r_26_sv2v_reg,
  scoreboard_r_25_sv2v_reg,scoreboard_r_24_sv2v_reg,scoreboard_r_23_sv2v_reg,
  scoreboard_r_22_sv2v_reg,scoreboard_r_21_sv2v_reg,scoreboard_r_20_sv2v_reg,
  scoreboard_r_19_sv2v_reg,scoreboard_r_18_sv2v_reg,scoreboard_r_17_sv2v_reg,scoreboard_r_16_sv2v_reg,
  scoreboard_r_15_sv2v_reg,scoreboard_r_14_sv2v_reg,scoreboard_r_13_sv2v_reg,
  scoreboard_r_12_sv2v_reg,scoreboard_r_11_sv2v_reg,scoreboard_r_10_sv2v_reg,
  scoreboard_r_9_sv2v_reg,scoreboard_r_8_sv2v_reg,scoreboard_r_7_sv2v_reg,
  scoreboard_r_6_sv2v_reg,scoreboard_r_5_sv2v_reg,scoreboard_r_4_sv2v_reg,scoreboard_r_3_sv2v_reg,
  scoreboard_r_2_sv2v_reg,scoreboard_r_1_sv2v_reg,scoreboard_r_0_sv2v_reg;
  assign scoreboard_r[31] = scoreboard_r_31_sv2v_reg;
  assign scoreboard_r[30] = scoreboard_r_30_sv2v_reg;
  assign scoreboard_r[29] = scoreboard_r_29_sv2v_reg;
  assign scoreboard_r[28] = scoreboard_r_28_sv2v_reg;
  assign scoreboard_r[27] = scoreboard_r_27_sv2v_reg;
  assign scoreboard_r[26] = scoreboard_r_26_sv2v_reg;
  assign scoreboard_r[25] = scoreboard_r_25_sv2v_reg;
  assign scoreboard_r[24] = scoreboard_r_24_sv2v_reg;
  assign scoreboard_r[23] = scoreboard_r_23_sv2v_reg;
  assign scoreboard_r[22] = scoreboard_r_22_sv2v_reg;
  assign scoreboard_r[21] = scoreboard_r_21_sv2v_reg;
  assign scoreboard_r[20] = scoreboard_r_20_sv2v_reg;
  assign scoreboard_r[19] = scoreboard_r_19_sv2v_reg;
  assign scoreboard_r[18] = scoreboard_r_18_sv2v_reg;
  assign scoreboard_r[17] = scoreboard_r_17_sv2v_reg;
  assign scoreboard_r[16] = scoreboard_r_16_sv2v_reg;
  assign scoreboard_r[15] = scoreboard_r_15_sv2v_reg;
  assign scoreboard_r[14] = scoreboard_r_14_sv2v_reg;
  assign scoreboard_r[13] = scoreboard_r_13_sv2v_reg;
  assign scoreboard_r[12] = scoreboard_r_12_sv2v_reg;
  assign scoreboard_r[11] = scoreboard_r_11_sv2v_reg;
  assign scoreboard_r[10] = scoreboard_r_10_sv2v_reg;
  assign scoreboard_r[9] = scoreboard_r_9_sv2v_reg;
  assign scoreboard_r[8] = scoreboard_r_8_sv2v_reg;
  assign scoreboard_r[7] = scoreboard_r_7_sv2v_reg;
  assign scoreboard_r[6] = scoreboard_r_6_sv2v_reg;
  assign scoreboard_r[5] = scoreboard_r_5_sv2v_reg;
  assign scoreboard_r[4] = scoreboard_r_4_sv2v_reg;
  assign scoreboard_r[3] = scoreboard_r_3_sv2v_reg;
  assign scoreboard_r[2] = scoreboard_r_2_sv2v_reg;
  assign scoreboard_r[1] = scoreboard_r_1_sv2v_reg;
  assign scoreboard_r[0] = scoreboard_r_0_sv2v_reg;

  bsg_transpose_width_p32_els_p1
  tranposer
  (
    .i(clear_by_port),
    .o(clear_by_port_t)
  );


  bsg_decode_with_v_num_out_p32
  \clr_dcode_v_0_.clear_decode_v 
  (
    .i(clear_id_i),
    .v_i(clear_i[0]),
    .o(clear_by_port)
  );


  bsg_decode_with_v_num_out_p32
  score_demux
  (
    .i(score_id_i),
    .v_i(_0_net_),
    .o(score_bits)
  );

  assign N65 = (N33)? scoreboard_r[0] : 
               (N35)? scoreboard_r[1] : 
               (N37)? scoreboard_r[2] : 
               (N39)? scoreboard_r[3] : 
               (N41)? scoreboard_r[4] : 
               (N43)? scoreboard_r[5] : 
               (N45)? scoreboard_r[6] : 
               (N47)? scoreboard_r[7] : 
               (N49)? scoreboard_r[8] : 
               (N51)? scoreboard_r[9] : 
               (N53)? scoreboard_r[10] : 
               (N55)? scoreboard_r[11] : 
               (N57)? scoreboard_r[12] : 
               (N59)? scoreboard_r[13] : 
               (N61)? scoreboard_r[14] : 
               (N63)? scoreboard_r[15] : 
               (N34)? scoreboard_r[16] : 
               (N36)? scoreboard_r[17] : 
               (N38)? scoreboard_r[18] : 
               (N40)? scoreboard_r[19] : 
               (N42)? scoreboard_r[20] : 
               (N44)? scoreboard_r[21] : 
               (N46)? scoreboard_r[22] : 
               (N48)? scoreboard_r[23] : 
               (N50)? scoreboard_r[24] : 
               (N52)? scoreboard_r[25] : 
               (N54)? scoreboard_r[26] : 
               (N56)? scoreboard_r[27] : 
               (N58)? scoreboard_r[28] : 
               (N60)? scoreboard_r[29] : 
               (N62)? scoreboard_r[30] : 
               (N64)? scoreboard_r[31] : 1'b0;
  assign N131 = (N99)? scoreboard_r[0] : 
                (N101)? scoreboard_r[1] : 
                (N103)? scoreboard_r[2] : 
                (N105)? scoreboard_r[3] : 
                (N107)? scoreboard_r[4] : 
                (N109)? scoreboard_r[5] : 
                (N111)? scoreboard_r[6] : 
                (N113)? scoreboard_r[7] : 
                (N115)? scoreboard_r[8] : 
                (N117)? scoreboard_r[9] : 
                (N119)? scoreboard_r[10] : 
                (N121)? scoreboard_r[11] : 
                (N123)? scoreboard_r[12] : 
                (N125)? scoreboard_r[13] : 
                (N127)? scoreboard_r[14] : 
                (N129)? scoreboard_r[15] : 
                (N100)? scoreboard_r[16] : 
                (N102)? scoreboard_r[17] : 
                (N104)? scoreboard_r[18] : 
                (N106)? scoreboard_r[19] : 
                (N108)? scoreboard_r[20] : 
                (N110)? scoreboard_r[21] : 
                (N112)? scoreboard_r[22] : 
                (N114)? scoreboard_r[23] : 
                (N116)? scoreboard_r[24] : 
                (N118)? scoreboard_r[25] : 
                (N120)? scoreboard_r[26] : 
                (N122)? scoreboard_r[27] : 
                (N124)? scoreboard_r[28] : 
                (N126)? scoreboard_r[29] : 
                (N128)? scoreboard_r[30] : 
                (N130)? scoreboard_r[31] : 1'b0;
  assign N197 = (N165)? scoreboard_r[0] : 
                (N167)? scoreboard_r[1] : 
                (N169)? scoreboard_r[2] : 
                (N171)? scoreboard_r[3] : 
                (N173)? scoreboard_r[4] : 
                (N175)? scoreboard_r[5] : 
                (N177)? scoreboard_r[6] : 
                (N179)? scoreboard_r[7] : 
                (N181)? scoreboard_r[8] : 
                (N183)? scoreboard_r[9] : 
                (N185)? scoreboard_r[10] : 
                (N187)? scoreboard_r[11] : 
                (N189)? scoreboard_r[12] : 
                (N191)? scoreboard_r[13] : 
                (N193)? scoreboard_r[14] : 
                (N195)? scoreboard_r[15] : 
                (N166)? scoreboard_r[16] : 
                (N168)? scoreboard_r[17] : 
                (N170)? scoreboard_r[18] : 
                (N172)? scoreboard_r[19] : 
                (N174)? scoreboard_r[20] : 
                (N176)? scoreboard_r[21] : 
                (N178)? scoreboard_r[22] : 
                (N180)? scoreboard_r[23] : 
                (N182)? scoreboard_r[24] : 
                (N184)? scoreboard_r[25] : 
                (N186)? scoreboard_r[26] : 
                (N188)? scoreboard_r[27] : 
                (N190)? scoreboard_r[28] : 
                (N192)? scoreboard_r[29] : 
                (N194)? scoreboard_r[30] : 
                (N196)? scoreboard_r[31] : 1'b0;
  assign N198 = clear_id_i == src_id_i[4:0];
  assign N199 = clear_id_i == src_id_i[9:5];
  assign N200 = clear_id_i == dest_id_i;

  bsg_transpose_width_p2_els_p1
  trans1
  (
    .i(rs_on_clear),
    .o(rs_on_clear_t)
  );

  assign N201 = src_id_i[4:0] == score_id_i;
  assign N202 = src_id_i[9:5] == score_id_i;
  assign N203 = dest_id_i == score_id_i;
  assign N204 = score_id_i[3] | score_id_i[4];
  assign N205 = score_id_i[2] | N204;
  assign N206 = score_id_i[1] | N205;
  assign N207 = score_id_i[0] | N206;
  assign _0_net_ = score_i & N207;
  assign N0 = ~src_id_i[0];
  assign N1 = ~src_id_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & src_id_i[1];
  assign N4 = src_id_i[0] & N1;
  assign N5 = src_id_i[0] & src_id_i[1];
  assign N6 = ~src_id_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & src_id_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & src_id_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & src_id_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & src_id_i[2];
  assign N15 = ~src_id_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & src_id_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & src_id_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & src_id_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & src_id_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & src_id_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & src_id_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & src_id_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & src_id_i[3];
  assign N32 = ~src_id_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & src_id_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & src_id_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & src_id_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & src_id_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & src_id_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & src_id_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & src_id_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & src_id_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & src_id_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & src_id_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & src_id_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & src_id_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & src_id_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & src_id_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & src_id_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & src_id_i[4];
  assign rs_depend_on_sb[0] = N65 & op_reads_rf_i[0];
  assign N66 = ~src_id_i[5];
  assign N67 = ~src_id_i[6];
  assign N68 = N66 & N67;
  assign N69 = N66 & src_id_i[6];
  assign N70 = src_id_i[5] & N67;
  assign N71 = src_id_i[5] & src_id_i[6];
  assign N72 = ~src_id_i[7];
  assign N73 = N68 & N72;
  assign N74 = N68 & src_id_i[7];
  assign N75 = N70 & N72;
  assign N76 = N70 & src_id_i[7];
  assign N77 = N69 & N72;
  assign N78 = N69 & src_id_i[7];
  assign N79 = N71 & N72;
  assign N80 = N71 & src_id_i[7];
  assign N81 = ~src_id_i[8];
  assign N82 = N73 & N81;
  assign N83 = N73 & src_id_i[8];
  assign N84 = N75 & N81;
  assign N85 = N75 & src_id_i[8];
  assign N86 = N77 & N81;
  assign N87 = N77 & src_id_i[8];
  assign N88 = N79 & N81;
  assign N89 = N79 & src_id_i[8];
  assign N90 = N74 & N81;
  assign N91 = N74 & src_id_i[8];
  assign N92 = N76 & N81;
  assign N93 = N76 & src_id_i[8];
  assign N94 = N78 & N81;
  assign N95 = N78 & src_id_i[8];
  assign N96 = N80 & N81;
  assign N97 = N80 & src_id_i[8];
  assign N98 = ~src_id_i[9];
  assign N99 = N82 & N98;
  assign N100 = N82 & src_id_i[9];
  assign N101 = N84 & N98;
  assign N102 = N84 & src_id_i[9];
  assign N103 = N86 & N98;
  assign N104 = N86 & src_id_i[9];
  assign N105 = N88 & N98;
  assign N106 = N88 & src_id_i[9];
  assign N107 = N90 & N98;
  assign N108 = N90 & src_id_i[9];
  assign N109 = N92 & N98;
  assign N110 = N92 & src_id_i[9];
  assign N111 = N94 & N98;
  assign N112 = N94 & src_id_i[9];
  assign N113 = N96 & N98;
  assign N114 = N96 & src_id_i[9];
  assign N115 = N83 & N98;
  assign N116 = N83 & src_id_i[9];
  assign N117 = N85 & N98;
  assign N118 = N85 & src_id_i[9];
  assign N119 = N87 & N98;
  assign N120 = N87 & src_id_i[9];
  assign N121 = N89 & N98;
  assign N122 = N89 & src_id_i[9];
  assign N123 = N91 & N98;
  assign N124 = N91 & src_id_i[9];
  assign N125 = N93 & N98;
  assign N126 = N93 & src_id_i[9];
  assign N127 = N95 & N98;
  assign N128 = N95 & src_id_i[9];
  assign N129 = N97 & N98;
  assign N130 = N97 & src_id_i[9];
  assign rs_depend_on_sb[1] = N131 & op_reads_rf_i[1];
  assign N132 = ~dest_id_i[0];
  assign N133 = ~dest_id_i[1];
  assign N134 = N132 & N133;
  assign N135 = N132 & dest_id_i[1];
  assign N136 = dest_id_i[0] & N133;
  assign N137 = dest_id_i[0] & dest_id_i[1];
  assign N138 = ~dest_id_i[2];
  assign N139 = N134 & N138;
  assign N140 = N134 & dest_id_i[2];
  assign N141 = N136 & N138;
  assign N142 = N136 & dest_id_i[2];
  assign N143 = N135 & N138;
  assign N144 = N135 & dest_id_i[2];
  assign N145 = N137 & N138;
  assign N146 = N137 & dest_id_i[2];
  assign N147 = ~dest_id_i[3];
  assign N148 = N139 & N147;
  assign N149 = N139 & dest_id_i[3];
  assign N150 = N141 & N147;
  assign N151 = N141 & dest_id_i[3];
  assign N152 = N143 & N147;
  assign N153 = N143 & dest_id_i[3];
  assign N154 = N145 & N147;
  assign N155 = N145 & dest_id_i[3];
  assign N156 = N140 & N147;
  assign N157 = N140 & dest_id_i[3];
  assign N158 = N142 & N147;
  assign N159 = N142 & dest_id_i[3];
  assign N160 = N144 & N147;
  assign N161 = N144 & dest_id_i[3];
  assign N162 = N146 & N147;
  assign N163 = N146 & dest_id_i[3];
  assign N164 = ~dest_id_i[4];
  assign N165 = N148 & N164;
  assign N166 = N148 & dest_id_i[4];
  assign N167 = N150 & N164;
  assign N168 = N150 & dest_id_i[4];
  assign N169 = N152 & N164;
  assign N170 = N152 & dest_id_i[4];
  assign N171 = N154 & N164;
  assign N172 = N154 & dest_id_i[4];
  assign N173 = N156 & N164;
  assign N174 = N156 & dest_id_i[4];
  assign N175 = N158 & N164;
  assign N176 = N158 & dest_id_i[4];
  assign N177 = N160 & N164;
  assign N178 = N160 & dest_id_i[4];
  assign N179 = N162 & N164;
  assign N180 = N162 & dest_id_i[4];
  assign N181 = N149 & N164;
  assign N182 = N149 & dest_id_i[4];
  assign N183 = N151 & N164;
  assign N184 = N151 & dest_id_i[4];
  assign N185 = N153 & N164;
  assign N186 = N153 & dest_id_i[4];
  assign N187 = N155 & N164;
  assign N188 = N155 & dest_id_i[4];
  assign N189 = N157 & N164;
  assign N190 = N157 & dest_id_i[4];
  assign N191 = N159 & N164;
  assign N192 = N159 & dest_id_i[4];
  assign N193 = N161 & N164;
  assign N194 = N161 & dest_id_i[4];
  assign N195 = N163 & N164;
  assign N196 = N163 & dest_id_i[4];
  assign rd_depend_on_sb = N197 & op_writes_rf_i;
  assign rs_on_clear[0] = clear_i[0] & N198;
  assign rs_on_clear[1] = clear_i[0] & N199;
  assign rd_on_clear[0] = clear_i[0] & N200;
  assign rs_depend_on_score[0] = N201 & op_reads_rf_i[0];
  assign rs_depend_on_score[1] = N202 & op_reads_rf_i[1];
  assign rd_depend_on_score = N203 & op_writes_rf_i;
  assign depend_on_sb = N212 | N214;
  assign N212 = N209 | N211;
  assign N209 = rd_depend_on_sb & N208;
  assign N208 = ~rd_on_clear[0];
  assign N211 = rs_depend_on_sb[1] & N210;
  assign N210 = ~rs_on_clear_t[1];
  assign N214 = rs_depend_on_sb[0] & N213;
  assign N213 = ~rs_on_clear_t[0];
  assign depend_on_score = N215 | rs_depend_on_score[0];
  assign N215 = rd_depend_on_score | rs_depend_on_score[1];
  assign dependency_o = depend_on_sb | N217;
  assign N217 = N216 & N207;
  assign N216 = depend_on_score & score_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      scoreboard_r_31_sv2v_reg <= 1'b0;
    end else if(score_bits[31]) begin
      scoreboard_r_31_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[31]) begin
      scoreboard_r_31_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_30_sv2v_reg <= 1'b0;
    end else if(score_bits[30]) begin
      scoreboard_r_30_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[30]) begin
      scoreboard_r_30_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_29_sv2v_reg <= 1'b0;
    end else if(score_bits[29]) begin
      scoreboard_r_29_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[29]) begin
      scoreboard_r_29_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_28_sv2v_reg <= 1'b0;
    end else if(score_bits[28]) begin
      scoreboard_r_28_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[28]) begin
      scoreboard_r_28_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_27_sv2v_reg <= 1'b0;
    end else if(score_bits[27]) begin
      scoreboard_r_27_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[27]) begin
      scoreboard_r_27_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_26_sv2v_reg <= 1'b0;
    end else if(score_bits[26]) begin
      scoreboard_r_26_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[26]) begin
      scoreboard_r_26_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_25_sv2v_reg <= 1'b0;
    end else if(score_bits[25]) begin
      scoreboard_r_25_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[25]) begin
      scoreboard_r_25_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_24_sv2v_reg <= 1'b0;
    end else if(score_bits[24]) begin
      scoreboard_r_24_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[24]) begin
      scoreboard_r_24_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_23_sv2v_reg <= 1'b0;
    end else if(score_bits[23]) begin
      scoreboard_r_23_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[23]) begin
      scoreboard_r_23_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_22_sv2v_reg <= 1'b0;
    end else if(score_bits[22]) begin
      scoreboard_r_22_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[22]) begin
      scoreboard_r_22_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_21_sv2v_reg <= 1'b0;
    end else if(score_bits[21]) begin
      scoreboard_r_21_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[21]) begin
      scoreboard_r_21_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_20_sv2v_reg <= 1'b0;
    end else if(score_bits[20]) begin
      scoreboard_r_20_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[20]) begin
      scoreboard_r_20_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_19_sv2v_reg <= 1'b0;
    end else if(score_bits[19]) begin
      scoreboard_r_19_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[19]) begin
      scoreboard_r_19_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_18_sv2v_reg <= 1'b0;
    end else if(score_bits[18]) begin
      scoreboard_r_18_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[18]) begin
      scoreboard_r_18_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_17_sv2v_reg <= 1'b0;
    end else if(score_bits[17]) begin
      scoreboard_r_17_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[17]) begin
      scoreboard_r_17_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_16_sv2v_reg <= 1'b0;
    end else if(score_bits[16]) begin
      scoreboard_r_16_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[16]) begin
      scoreboard_r_16_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_15_sv2v_reg <= 1'b0;
    end else if(score_bits[15]) begin
      scoreboard_r_15_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[15]) begin
      scoreboard_r_15_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_14_sv2v_reg <= 1'b0;
    end else if(score_bits[14]) begin
      scoreboard_r_14_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[14]) begin
      scoreboard_r_14_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_13_sv2v_reg <= 1'b0;
    end else if(score_bits[13]) begin
      scoreboard_r_13_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[13]) begin
      scoreboard_r_13_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_12_sv2v_reg <= 1'b0;
    end else if(score_bits[12]) begin
      scoreboard_r_12_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[12]) begin
      scoreboard_r_12_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_11_sv2v_reg <= 1'b0;
    end else if(score_bits[11]) begin
      scoreboard_r_11_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[11]) begin
      scoreboard_r_11_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_10_sv2v_reg <= 1'b0;
    end else if(score_bits[10]) begin
      scoreboard_r_10_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[10]) begin
      scoreboard_r_10_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_9_sv2v_reg <= 1'b0;
    end else if(score_bits[9]) begin
      scoreboard_r_9_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[9]) begin
      scoreboard_r_9_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_8_sv2v_reg <= 1'b0;
    end else if(score_bits[8]) begin
      scoreboard_r_8_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[8]) begin
      scoreboard_r_8_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_7_sv2v_reg <= 1'b0;
    end else if(score_bits[7]) begin
      scoreboard_r_7_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[7]) begin
      scoreboard_r_7_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_6_sv2v_reg <= 1'b0;
    end else if(score_bits[6]) begin
      scoreboard_r_6_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[6]) begin
      scoreboard_r_6_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_5_sv2v_reg <= 1'b0;
    end else if(score_bits[5]) begin
      scoreboard_r_5_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[5]) begin
      scoreboard_r_5_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_4_sv2v_reg <= 1'b0;
    end else if(score_bits[4]) begin
      scoreboard_r_4_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[4]) begin
      scoreboard_r_4_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_3_sv2v_reg <= 1'b0;
    end else if(score_bits[3]) begin
      scoreboard_r_3_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[3]) begin
      scoreboard_r_3_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_2_sv2v_reg <= 1'b0;
    end else if(score_bits[2]) begin
      scoreboard_r_2_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[2]) begin
      scoreboard_r_2_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_1_sv2v_reg <= 1'b0;
    end else if(score_bits[1]) begin
      scoreboard_r_1_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[1]) begin
      scoreboard_r_1_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_0_sv2v_reg <= 1'b0;
    end else if(score_bits[0]) begin
      scoreboard_r_0_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[0]) begin
      scoreboard_r_0_sv2v_reg <= 1'b0;
    end 
  end


endmodule



module regfile_synth_width_p33_els_p32_num_rs_p3_x0_tied_to_zero_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [4:0] w_addr_i;
  input [32:0] w_data_i;
  input [2:0] r_v_i;
  input [14:0] r_addr_i;
  output [98:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  wire [98:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286;
  wire [14:0] r_addr_r;
  wire [1055:0] \xnz.mem_r ;
  reg r_addr_r_14_sv2v_reg,r_addr_r_13_sv2v_reg,r_addr_r_12_sv2v_reg,
  r_addr_r_11_sv2v_reg,r_addr_r_10_sv2v_reg,r_addr_r_9_sv2v_reg,r_addr_r_8_sv2v_reg,
  r_addr_r_7_sv2v_reg,r_addr_r_6_sv2v_reg,r_addr_r_5_sv2v_reg,r_addr_r_4_sv2v_reg,
  r_addr_r_3_sv2v_reg,r_addr_r_2_sv2v_reg,r_addr_r_1_sv2v_reg,r_addr_r_0_sv2v_reg,
  \xnz.mem_r_1055_sv2v_reg ,\xnz.mem_r_1054_sv2v_reg ,\xnz.mem_r_1053_sv2v_reg ,
  \xnz.mem_r_1052_sv2v_reg ,\xnz.mem_r_1051_sv2v_reg ,\xnz.mem_r_1050_sv2v_reg ,
  \xnz.mem_r_1049_sv2v_reg ,\xnz.mem_r_1048_sv2v_reg ,\xnz.mem_r_1047_sv2v_reg ,
  \xnz.mem_r_1046_sv2v_reg ,\xnz.mem_r_1045_sv2v_reg ,\xnz.mem_r_1044_sv2v_reg ,
  \xnz.mem_r_1043_sv2v_reg ,\xnz.mem_r_1042_sv2v_reg ,\xnz.mem_r_1041_sv2v_reg ,
  \xnz.mem_r_1040_sv2v_reg ,\xnz.mem_r_1039_sv2v_reg ,\xnz.mem_r_1038_sv2v_reg ,\xnz.mem_r_1037_sv2v_reg ,
  \xnz.mem_r_1036_sv2v_reg ,\xnz.mem_r_1035_sv2v_reg ,\xnz.mem_r_1034_sv2v_reg ,
  \xnz.mem_r_1033_sv2v_reg ,\xnz.mem_r_1032_sv2v_reg ,\xnz.mem_r_1031_sv2v_reg ,
  \xnz.mem_r_1030_sv2v_reg ,\xnz.mem_r_1029_sv2v_reg ,\xnz.mem_r_1028_sv2v_reg ,
  \xnz.mem_r_1027_sv2v_reg ,\xnz.mem_r_1026_sv2v_reg ,\xnz.mem_r_1025_sv2v_reg ,
  \xnz.mem_r_1024_sv2v_reg ,\xnz.mem_r_1023_sv2v_reg ,\xnz.mem_r_1022_sv2v_reg ,
  \xnz.mem_r_1021_sv2v_reg ,\xnz.mem_r_1020_sv2v_reg ,\xnz.mem_r_1019_sv2v_reg ,
  \xnz.mem_r_1018_sv2v_reg ,\xnz.mem_r_1017_sv2v_reg ,\xnz.mem_r_1016_sv2v_reg ,
  \xnz.mem_r_1015_sv2v_reg ,\xnz.mem_r_1014_sv2v_reg ,\xnz.mem_r_1013_sv2v_reg ,
  \xnz.mem_r_1012_sv2v_reg ,\xnz.mem_r_1011_sv2v_reg ,\xnz.mem_r_1010_sv2v_reg ,
  \xnz.mem_r_1009_sv2v_reg ,\xnz.mem_r_1008_sv2v_reg ,\xnz.mem_r_1007_sv2v_reg ,
  \xnz.mem_r_1006_sv2v_reg ,\xnz.mem_r_1005_sv2v_reg ,\xnz.mem_r_1004_sv2v_reg ,
  \xnz.mem_r_1003_sv2v_reg ,\xnz.mem_r_1002_sv2v_reg ,\xnz.mem_r_1001_sv2v_reg ,
  \xnz.mem_r_1000_sv2v_reg ,\xnz.mem_r_999_sv2v_reg ,\xnz.mem_r_998_sv2v_reg ,\xnz.mem_r_997_sv2v_reg ,
  \xnz.mem_r_996_sv2v_reg ,\xnz.mem_r_995_sv2v_reg ,\xnz.mem_r_994_sv2v_reg ,
  \xnz.mem_r_993_sv2v_reg ,\xnz.mem_r_992_sv2v_reg ,\xnz.mem_r_991_sv2v_reg ,
  \xnz.mem_r_990_sv2v_reg ,\xnz.mem_r_989_sv2v_reg ,\xnz.mem_r_988_sv2v_reg ,
  \xnz.mem_r_987_sv2v_reg ,\xnz.mem_r_986_sv2v_reg ,\xnz.mem_r_985_sv2v_reg ,
  \xnz.mem_r_984_sv2v_reg ,\xnz.mem_r_983_sv2v_reg ,\xnz.mem_r_982_sv2v_reg ,\xnz.mem_r_981_sv2v_reg ,
  \xnz.mem_r_980_sv2v_reg ,\xnz.mem_r_979_sv2v_reg ,\xnz.mem_r_978_sv2v_reg ,
  \xnz.mem_r_977_sv2v_reg ,\xnz.mem_r_976_sv2v_reg ,\xnz.mem_r_975_sv2v_reg ,
  \xnz.mem_r_974_sv2v_reg ,\xnz.mem_r_973_sv2v_reg ,\xnz.mem_r_972_sv2v_reg ,
  \xnz.mem_r_971_sv2v_reg ,\xnz.mem_r_970_sv2v_reg ,\xnz.mem_r_969_sv2v_reg ,
  \xnz.mem_r_968_sv2v_reg ,\xnz.mem_r_967_sv2v_reg ,\xnz.mem_r_966_sv2v_reg ,\xnz.mem_r_965_sv2v_reg ,
  \xnz.mem_r_964_sv2v_reg ,\xnz.mem_r_963_sv2v_reg ,\xnz.mem_r_962_sv2v_reg ,
  \xnz.mem_r_961_sv2v_reg ,\xnz.mem_r_960_sv2v_reg ,\xnz.mem_r_959_sv2v_reg ,
  \xnz.mem_r_958_sv2v_reg ,\xnz.mem_r_957_sv2v_reg ,\xnz.mem_r_956_sv2v_reg ,
  \xnz.mem_r_955_sv2v_reg ,\xnz.mem_r_954_sv2v_reg ,\xnz.mem_r_953_sv2v_reg ,
  \xnz.mem_r_952_sv2v_reg ,\xnz.mem_r_951_sv2v_reg ,\xnz.mem_r_950_sv2v_reg ,\xnz.mem_r_949_sv2v_reg ,
  \xnz.mem_r_948_sv2v_reg ,\xnz.mem_r_947_sv2v_reg ,\xnz.mem_r_946_sv2v_reg ,
  \xnz.mem_r_945_sv2v_reg ,\xnz.mem_r_944_sv2v_reg ,\xnz.mem_r_943_sv2v_reg ,
  \xnz.mem_r_942_sv2v_reg ,\xnz.mem_r_941_sv2v_reg ,\xnz.mem_r_940_sv2v_reg ,
  \xnz.mem_r_939_sv2v_reg ,\xnz.mem_r_938_sv2v_reg ,\xnz.mem_r_937_sv2v_reg ,
  \xnz.mem_r_936_sv2v_reg ,\xnz.mem_r_935_sv2v_reg ,\xnz.mem_r_934_sv2v_reg ,\xnz.mem_r_933_sv2v_reg ,
  \xnz.mem_r_932_sv2v_reg ,\xnz.mem_r_931_sv2v_reg ,\xnz.mem_r_930_sv2v_reg ,
  \xnz.mem_r_929_sv2v_reg ,\xnz.mem_r_928_sv2v_reg ,\xnz.mem_r_927_sv2v_reg ,
  \xnz.mem_r_926_sv2v_reg ,\xnz.mem_r_925_sv2v_reg ,\xnz.mem_r_924_sv2v_reg ,
  \xnz.mem_r_923_sv2v_reg ,\xnz.mem_r_922_sv2v_reg ,\xnz.mem_r_921_sv2v_reg ,
  \xnz.mem_r_920_sv2v_reg ,\xnz.mem_r_919_sv2v_reg ,\xnz.mem_r_918_sv2v_reg ,\xnz.mem_r_917_sv2v_reg ,
  \xnz.mem_r_916_sv2v_reg ,\xnz.mem_r_915_sv2v_reg ,\xnz.mem_r_914_sv2v_reg ,
  \xnz.mem_r_913_sv2v_reg ,\xnz.mem_r_912_sv2v_reg ,\xnz.mem_r_911_sv2v_reg ,
  \xnz.mem_r_910_sv2v_reg ,\xnz.mem_r_909_sv2v_reg ,\xnz.mem_r_908_sv2v_reg ,
  \xnz.mem_r_907_sv2v_reg ,\xnz.mem_r_906_sv2v_reg ,\xnz.mem_r_905_sv2v_reg ,
  \xnz.mem_r_904_sv2v_reg ,\xnz.mem_r_903_sv2v_reg ,\xnz.mem_r_902_sv2v_reg ,\xnz.mem_r_901_sv2v_reg ,
  \xnz.mem_r_900_sv2v_reg ,\xnz.mem_r_899_sv2v_reg ,\xnz.mem_r_898_sv2v_reg ,
  \xnz.mem_r_897_sv2v_reg ,\xnz.mem_r_896_sv2v_reg ,\xnz.mem_r_895_sv2v_reg ,
  \xnz.mem_r_894_sv2v_reg ,\xnz.mem_r_893_sv2v_reg ,\xnz.mem_r_892_sv2v_reg ,
  \xnz.mem_r_891_sv2v_reg ,\xnz.mem_r_890_sv2v_reg ,\xnz.mem_r_889_sv2v_reg ,
  \xnz.mem_r_888_sv2v_reg ,\xnz.mem_r_887_sv2v_reg ,\xnz.mem_r_886_sv2v_reg ,\xnz.mem_r_885_sv2v_reg ,
  \xnz.mem_r_884_sv2v_reg ,\xnz.mem_r_883_sv2v_reg ,\xnz.mem_r_882_sv2v_reg ,
  \xnz.mem_r_881_sv2v_reg ,\xnz.mem_r_880_sv2v_reg ,\xnz.mem_r_879_sv2v_reg ,
  \xnz.mem_r_878_sv2v_reg ,\xnz.mem_r_877_sv2v_reg ,\xnz.mem_r_876_sv2v_reg ,
  \xnz.mem_r_875_sv2v_reg ,\xnz.mem_r_874_sv2v_reg ,\xnz.mem_r_873_sv2v_reg ,
  \xnz.mem_r_872_sv2v_reg ,\xnz.mem_r_871_sv2v_reg ,\xnz.mem_r_870_sv2v_reg ,\xnz.mem_r_869_sv2v_reg ,
  \xnz.mem_r_868_sv2v_reg ,\xnz.mem_r_867_sv2v_reg ,\xnz.mem_r_866_sv2v_reg ,
  \xnz.mem_r_865_sv2v_reg ,\xnz.mem_r_864_sv2v_reg ,\xnz.mem_r_863_sv2v_reg ,
  \xnz.mem_r_862_sv2v_reg ,\xnz.mem_r_861_sv2v_reg ,\xnz.mem_r_860_sv2v_reg ,
  \xnz.mem_r_859_sv2v_reg ,\xnz.mem_r_858_sv2v_reg ,\xnz.mem_r_857_sv2v_reg ,
  \xnz.mem_r_856_sv2v_reg ,\xnz.mem_r_855_sv2v_reg ,\xnz.mem_r_854_sv2v_reg ,\xnz.mem_r_853_sv2v_reg ,
  \xnz.mem_r_852_sv2v_reg ,\xnz.mem_r_851_sv2v_reg ,\xnz.mem_r_850_sv2v_reg ,
  \xnz.mem_r_849_sv2v_reg ,\xnz.mem_r_848_sv2v_reg ,\xnz.mem_r_847_sv2v_reg ,
  \xnz.mem_r_846_sv2v_reg ,\xnz.mem_r_845_sv2v_reg ,\xnz.mem_r_844_sv2v_reg ,
  \xnz.mem_r_843_sv2v_reg ,\xnz.mem_r_842_sv2v_reg ,\xnz.mem_r_841_sv2v_reg ,
  \xnz.mem_r_840_sv2v_reg ,\xnz.mem_r_839_sv2v_reg ,\xnz.mem_r_838_sv2v_reg ,\xnz.mem_r_837_sv2v_reg ,
  \xnz.mem_r_836_sv2v_reg ,\xnz.mem_r_835_sv2v_reg ,\xnz.mem_r_834_sv2v_reg ,
  \xnz.mem_r_833_sv2v_reg ,\xnz.mem_r_832_sv2v_reg ,\xnz.mem_r_831_sv2v_reg ,
  \xnz.mem_r_830_sv2v_reg ,\xnz.mem_r_829_sv2v_reg ,\xnz.mem_r_828_sv2v_reg ,
  \xnz.mem_r_827_sv2v_reg ,\xnz.mem_r_826_sv2v_reg ,\xnz.mem_r_825_sv2v_reg ,
  \xnz.mem_r_824_sv2v_reg ,\xnz.mem_r_823_sv2v_reg ,\xnz.mem_r_822_sv2v_reg ,\xnz.mem_r_821_sv2v_reg ,
  \xnz.mem_r_820_sv2v_reg ,\xnz.mem_r_819_sv2v_reg ,\xnz.mem_r_818_sv2v_reg ,
  \xnz.mem_r_817_sv2v_reg ,\xnz.mem_r_816_sv2v_reg ,\xnz.mem_r_815_sv2v_reg ,
  \xnz.mem_r_814_sv2v_reg ,\xnz.mem_r_813_sv2v_reg ,\xnz.mem_r_812_sv2v_reg ,
  \xnz.mem_r_811_sv2v_reg ,\xnz.mem_r_810_sv2v_reg ,\xnz.mem_r_809_sv2v_reg ,
  \xnz.mem_r_808_sv2v_reg ,\xnz.mem_r_807_sv2v_reg ,\xnz.mem_r_806_sv2v_reg ,\xnz.mem_r_805_sv2v_reg ,
  \xnz.mem_r_804_sv2v_reg ,\xnz.mem_r_803_sv2v_reg ,\xnz.mem_r_802_sv2v_reg ,
  \xnz.mem_r_801_sv2v_reg ,\xnz.mem_r_800_sv2v_reg ,\xnz.mem_r_799_sv2v_reg ,
  \xnz.mem_r_798_sv2v_reg ,\xnz.mem_r_797_sv2v_reg ,\xnz.mem_r_796_sv2v_reg ,
  \xnz.mem_r_795_sv2v_reg ,\xnz.mem_r_794_sv2v_reg ,\xnz.mem_r_793_sv2v_reg ,
  \xnz.mem_r_792_sv2v_reg ,\xnz.mem_r_791_sv2v_reg ,\xnz.mem_r_790_sv2v_reg ,\xnz.mem_r_789_sv2v_reg ,
  \xnz.mem_r_788_sv2v_reg ,\xnz.mem_r_787_sv2v_reg ,\xnz.mem_r_786_sv2v_reg ,
  \xnz.mem_r_785_sv2v_reg ,\xnz.mem_r_784_sv2v_reg ,\xnz.mem_r_783_sv2v_reg ,
  \xnz.mem_r_782_sv2v_reg ,\xnz.mem_r_781_sv2v_reg ,\xnz.mem_r_780_sv2v_reg ,
  \xnz.mem_r_779_sv2v_reg ,\xnz.mem_r_778_sv2v_reg ,\xnz.mem_r_777_sv2v_reg ,
  \xnz.mem_r_776_sv2v_reg ,\xnz.mem_r_775_sv2v_reg ,\xnz.mem_r_774_sv2v_reg ,\xnz.mem_r_773_sv2v_reg ,
  \xnz.mem_r_772_sv2v_reg ,\xnz.mem_r_771_sv2v_reg ,\xnz.mem_r_770_sv2v_reg ,
  \xnz.mem_r_769_sv2v_reg ,\xnz.mem_r_768_sv2v_reg ,\xnz.mem_r_767_sv2v_reg ,
  \xnz.mem_r_766_sv2v_reg ,\xnz.mem_r_765_sv2v_reg ,\xnz.mem_r_764_sv2v_reg ,
  \xnz.mem_r_763_sv2v_reg ,\xnz.mem_r_762_sv2v_reg ,\xnz.mem_r_761_sv2v_reg ,
  \xnz.mem_r_760_sv2v_reg ,\xnz.mem_r_759_sv2v_reg ,\xnz.mem_r_758_sv2v_reg ,\xnz.mem_r_757_sv2v_reg ,
  \xnz.mem_r_756_sv2v_reg ,\xnz.mem_r_755_sv2v_reg ,\xnz.mem_r_754_sv2v_reg ,
  \xnz.mem_r_753_sv2v_reg ,\xnz.mem_r_752_sv2v_reg ,\xnz.mem_r_751_sv2v_reg ,
  \xnz.mem_r_750_sv2v_reg ,\xnz.mem_r_749_sv2v_reg ,\xnz.mem_r_748_sv2v_reg ,
  \xnz.mem_r_747_sv2v_reg ,\xnz.mem_r_746_sv2v_reg ,\xnz.mem_r_745_sv2v_reg ,
  \xnz.mem_r_744_sv2v_reg ,\xnz.mem_r_743_sv2v_reg ,\xnz.mem_r_742_sv2v_reg ,\xnz.mem_r_741_sv2v_reg ,
  \xnz.mem_r_740_sv2v_reg ,\xnz.mem_r_739_sv2v_reg ,\xnz.mem_r_738_sv2v_reg ,
  \xnz.mem_r_737_sv2v_reg ,\xnz.mem_r_736_sv2v_reg ,\xnz.mem_r_735_sv2v_reg ,
  \xnz.mem_r_734_sv2v_reg ,\xnz.mem_r_733_sv2v_reg ,\xnz.mem_r_732_sv2v_reg ,
  \xnz.mem_r_731_sv2v_reg ,\xnz.mem_r_730_sv2v_reg ,\xnz.mem_r_729_sv2v_reg ,
  \xnz.mem_r_728_sv2v_reg ,\xnz.mem_r_727_sv2v_reg ,\xnz.mem_r_726_sv2v_reg ,\xnz.mem_r_725_sv2v_reg ,
  \xnz.mem_r_724_sv2v_reg ,\xnz.mem_r_723_sv2v_reg ,\xnz.mem_r_722_sv2v_reg ,
  \xnz.mem_r_721_sv2v_reg ,\xnz.mem_r_720_sv2v_reg ,\xnz.mem_r_719_sv2v_reg ,
  \xnz.mem_r_718_sv2v_reg ,\xnz.mem_r_717_sv2v_reg ,\xnz.mem_r_716_sv2v_reg ,
  \xnz.mem_r_715_sv2v_reg ,\xnz.mem_r_714_sv2v_reg ,\xnz.mem_r_713_sv2v_reg ,
  \xnz.mem_r_712_sv2v_reg ,\xnz.mem_r_711_sv2v_reg ,\xnz.mem_r_710_sv2v_reg ,\xnz.mem_r_709_sv2v_reg ,
  \xnz.mem_r_708_sv2v_reg ,\xnz.mem_r_707_sv2v_reg ,\xnz.mem_r_706_sv2v_reg ,
  \xnz.mem_r_705_sv2v_reg ,\xnz.mem_r_704_sv2v_reg ,\xnz.mem_r_703_sv2v_reg ,
  \xnz.mem_r_702_sv2v_reg ,\xnz.mem_r_701_sv2v_reg ,\xnz.mem_r_700_sv2v_reg ,
  \xnz.mem_r_699_sv2v_reg ,\xnz.mem_r_698_sv2v_reg ,\xnz.mem_r_697_sv2v_reg ,
  \xnz.mem_r_696_sv2v_reg ,\xnz.mem_r_695_sv2v_reg ,\xnz.mem_r_694_sv2v_reg ,\xnz.mem_r_693_sv2v_reg ,
  \xnz.mem_r_692_sv2v_reg ,\xnz.mem_r_691_sv2v_reg ,\xnz.mem_r_690_sv2v_reg ,
  \xnz.mem_r_689_sv2v_reg ,\xnz.mem_r_688_sv2v_reg ,\xnz.mem_r_687_sv2v_reg ,
  \xnz.mem_r_686_sv2v_reg ,\xnz.mem_r_685_sv2v_reg ,\xnz.mem_r_684_sv2v_reg ,
  \xnz.mem_r_683_sv2v_reg ,\xnz.mem_r_682_sv2v_reg ,\xnz.mem_r_681_sv2v_reg ,
  \xnz.mem_r_680_sv2v_reg ,\xnz.mem_r_679_sv2v_reg ,\xnz.mem_r_678_sv2v_reg ,\xnz.mem_r_677_sv2v_reg ,
  \xnz.mem_r_676_sv2v_reg ,\xnz.mem_r_675_sv2v_reg ,\xnz.mem_r_674_sv2v_reg ,
  \xnz.mem_r_673_sv2v_reg ,\xnz.mem_r_672_sv2v_reg ,\xnz.mem_r_671_sv2v_reg ,
  \xnz.mem_r_670_sv2v_reg ,\xnz.mem_r_669_sv2v_reg ,\xnz.mem_r_668_sv2v_reg ,
  \xnz.mem_r_667_sv2v_reg ,\xnz.mem_r_666_sv2v_reg ,\xnz.mem_r_665_sv2v_reg ,
  \xnz.mem_r_664_sv2v_reg ,\xnz.mem_r_663_sv2v_reg ,\xnz.mem_r_662_sv2v_reg ,\xnz.mem_r_661_sv2v_reg ,
  \xnz.mem_r_660_sv2v_reg ,\xnz.mem_r_659_sv2v_reg ,\xnz.mem_r_658_sv2v_reg ,
  \xnz.mem_r_657_sv2v_reg ,\xnz.mem_r_656_sv2v_reg ,\xnz.mem_r_655_sv2v_reg ,
  \xnz.mem_r_654_sv2v_reg ,\xnz.mem_r_653_sv2v_reg ,\xnz.mem_r_652_sv2v_reg ,
  \xnz.mem_r_651_sv2v_reg ,\xnz.mem_r_650_sv2v_reg ,\xnz.mem_r_649_sv2v_reg ,
  \xnz.mem_r_648_sv2v_reg ,\xnz.mem_r_647_sv2v_reg ,\xnz.mem_r_646_sv2v_reg ,\xnz.mem_r_645_sv2v_reg ,
  \xnz.mem_r_644_sv2v_reg ,\xnz.mem_r_643_sv2v_reg ,\xnz.mem_r_642_sv2v_reg ,
  \xnz.mem_r_641_sv2v_reg ,\xnz.mem_r_640_sv2v_reg ,\xnz.mem_r_639_sv2v_reg ,
  \xnz.mem_r_638_sv2v_reg ,\xnz.mem_r_637_sv2v_reg ,\xnz.mem_r_636_sv2v_reg ,
  \xnz.mem_r_635_sv2v_reg ,\xnz.mem_r_634_sv2v_reg ,\xnz.mem_r_633_sv2v_reg ,
  \xnz.mem_r_632_sv2v_reg ,\xnz.mem_r_631_sv2v_reg ,\xnz.mem_r_630_sv2v_reg ,\xnz.mem_r_629_sv2v_reg ,
  \xnz.mem_r_628_sv2v_reg ,\xnz.mem_r_627_sv2v_reg ,\xnz.mem_r_626_sv2v_reg ,
  \xnz.mem_r_625_sv2v_reg ,\xnz.mem_r_624_sv2v_reg ,\xnz.mem_r_623_sv2v_reg ,
  \xnz.mem_r_622_sv2v_reg ,\xnz.mem_r_621_sv2v_reg ,\xnz.mem_r_620_sv2v_reg ,
  \xnz.mem_r_619_sv2v_reg ,\xnz.mem_r_618_sv2v_reg ,\xnz.mem_r_617_sv2v_reg ,
  \xnz.mem_r_616_sv2v_reg ,\xnz.mem_r_615_sv2v_reg ,\xnz.mem_r_614_sv2v_reg ,\xnz.mem_r_613_sv2v_reg ,
  \xnz.mem_r_612_sv2v_reg ,\xnz.mem_r_611_sv2v_reg ,\xnz.mem_r_610_sv2v_reg ,
  \xnz.mem_r_609_sv2v_reg ,\xnz.mem_r_608_sv2v_reg ,\xnz.mem_r_607_sv2v_reg ,
  \xnz.mem_r_606_sv2v_reg ,\xnz.mem_r_605_sv2v_reg ,\xnz.mem_r_604_sv2v_reg ,
  \xnz.mem_r_603_sv2v_reg ,\xnz.mem_r_602_sv2v_reg ,\xnz.mem_r_601_sv2v_reg ,
  \xnz.mem_r_600_sv2v_reg ,\xnz.mem_r_599_sv2v_reg ,\xnz.mem_r_598_sv2v_reg ,\xnz.mem_r_597_sv2v_reg ,
  \xnz.mem_r_596_sv2v_reg ,\xnz.mem_r_595_sv2v_reg ,\xnz.mem_r_594_sv2v_reg ,
  \xnz.mem_r_593_sv2v_reg ,\xnz.mem_r_592_sv2v_reg ,\xnz.mem_r_591_sv2v_reg ,
  \xnz.mem_r_590_sv2v_reg ,\xnz.mem_r_589_sv2v_reg ,\xnz.mem_r_588_sv2v_reg ,
  \xnz.mem_r_587_sv2v_reg ,\xnz.mem_r_586_sv2v_reg ,\xnz.mem_r_585_sv2v_reg ,
  \xnz.mem_r_584_sv2v_reg ,\xnz.mem_r_583_sv2v_reg ,\xnz.mem_r_582_sv2v_reg ,\xnz.mem_r_581_sv2v_reg ,
  \xnz.mem_r_580_sv2v_reg ,\xnz.mem_r_579_sv2v_reg ,\xnz.mem_r_578_sv2v_reg ,
  \xnz.mem_r_577_sv2v_reg ,\xnz.mem_r_576_sv2v_reg ,\xnz.mem_r_575_sv2v_reg ,
  \xnz.mem_r_574_sv2v_reg ,\xnz.mem_r_573_sv2v_reg ,\xnz.mem_r_572_sv2v_reg ,
  \xnz.mem_r_571_sv2v_reg ,\xnz.mem_r_570_sv2v_reg ,\xnz.mem_r_569_sv2v_reg ,
  \xnz.mem_r_568_sv2v_reg ,\xnz.mem_r_567_sv2v_reg ,\xnz.mem_r_566_sv2v_reg ,\xnz.mem_r_565_sv2v_reg ,
  \xnz.mem_r_564_sv2v_reg ,\xnz.mem_r_563_sv2v_reg ,\xnz.mem_r_562_sv2v_reg ,
  \xnz.mem_r_561_sv2v_reg ,\xnz.mem_r_560_sv2v_reg ,\xnz.mem_r_559_sv2v_reg ,
  \xnz.mem_r_558_sv2v_reg ,\xnz.mem_r_557_sv2v_reg ,\xnz.mem_r_556_sv2v_reg ,
  \xnz.mem_r_555_sv2v_reg ,\xnz.mem_r_554_sv2v_reg ,\xnz.mem_r_553_sv2v_reg ,
  \xnz.mem_r_552_sv2v_reg ,\xnz.mem_r_551_sv2v_reg ,\xnz.mem_r_550_sv2v_reg ,\xnz.mem_r_549_sv2v_reg ,
  \xnz.mem_r_548_sv2v_reg ,\xnz.mem_r_547_sv2v_reg ,\xnz.mem_r_546_sv2v_reg ,
  \xnz.mem_r_545_sv2v_reg ,\xnz.mem_r_544_sv2v_reg ,\xnz.mem_r_543_sv2v_reg ,
  \xnz.mem_r_542_sv2v_reg ,\xnz.mem_r_541_sv2v_reg ,\xnz.mem_r_540_sv2v_reg ,
  \xnz.mem_r_539_sv2v_reg ,\xnz.mem_r_538_sv2v_reg ,\xnz.mem_r_537_sv2v_reg ,
  \xnz.mem_r_536_sv2v_reg ,\xnz.mem_r_535_sv2v_reg ,\xnz.mem_r_534_sv2v_reg ,\xnz.mem_r_533_sv2v_reg ,
  \xnz.mem_r_532_sv2v_reg ,\xnz.mem_r_531_sv2v_reg ,\xnz.mem_r_530_sv2v_reg ,
  \xnz.mem_r_529_sv2v_reg ,\xnz.mem_r_528_sv2v_reg ,\xnz.mem_r_527_sv2v_reg ,
  \xnz.mem_r_526_sv2v_reg ,\xnz.mem_r_525_sv2v_reg ,\xnz.mem_r_524_sv2v_reg ,
  \xnz.mem_r_523_sv2v_reg ,\xnz.mem_r_522_sv2v_reg ,\xnz.mem_r_521_sv2v_reg ,
  \xnz.mem_r_520_sv2v_reg ,\xnz.mem_r_519_sv2v_reg ,\xnz.mem_r_518_sv2v_reg ,\xnz.mem_r_517_sv2v_reg ,
  \xnz.mem_r_516_sv2v_reg ,\xnz.mem_r_515_sv2v_reg ,\xnz.mem_r_514_sv2v_reg ,
  \xnz.mem_r_513_sv2v_reg ,\xnz.mem_r_512_sv2v_reg ,\xnz.mem_r_511_sv2v_reg ,
  \xnz.mem_r_510_sv2v_reg ,\xnz.mem_r_509_sv2v_reg ,\xnz.mem_r_508_sv2v_reg ,
  \xnz.mem_r_507_sv2v_reg ,\xnz.mem_r_506_sv2v_reg ,\xnz.mem_r_505_sv2v_reg ,
  \xnz.mem_r_504_sv2v_reg ,\xnz.mem_r_503_sv2v_reg ,\xnz.mem_r_502_sv2v_reg ,\xnz.mem_r_501_sv2v_reg ,
  \xnz.mem_r_500_sv2v_reg ,\xnz.mem_r_499_sv2v_reg ,\xnz.mem_r_498_sv2v_reg ,
  \xnz.mem_r_497_sv2v_reg ,\xnz.mem_r_496_sv2v_reg ,\xnz.mem_r_495_sv2v_reg ,
  \xnz.mem_r_494_sv2v_reg ,\xnz.mem_r_493_sv2v_reg ,\xnz.mem_r_492_sv2v_reg ,
  \xnz.mem_r_491_sv2v_reg ,\xnz.mem_r_490_sv2v_reg ,\xnz.mem_r_489_sv2v_reg ,
  \xnz.mem_r_488_sv2v_reg ,\xnz.mem_r_487_sv2v_reg ,\xnz.mem_r_486_sv2v_reg ,\xnz.mem_r_485_sv2v_reg ,
  \xnz.mem_r_484_sv2v_reg ,\xnz.mem_r_483_sv2v_reg ,\xnz.mem_r_482_sv2v_reg ,
  \xnz.mem_r_481_sv2v_reg ,\xnz.mem_r_480_sv2v_reg ,\xnz.mem_r_479_sv2v_reg ,
  \xnz.mem_r_478_sv2v_reg ,\xnz.mem_r_477_sv2v_reg ,\xnz.mem_r_476_sv2v_reg ,
  \xnz.mem_r_475_sv2v_reg ,\xnz.mem_r_474_sv2v_reg ,\xnz.mem_r_473_sv2v_reg ,
  \xnz.mem_r_472_sv2v_reg ,\xnz.mem_r_471_sv2v_reg ,\xnz.mem_r_470_sv2v_reg ,\xnz.mem_r_469_sv2v_reg ,
  \xnz.mem_r_468_sv2v_reg ,\xnz.mem_r_467_sv2v_reg ,\xnz.mem_r_466_sv2v_reg ,
  \xnz.mem_r_465_sv2v_reg ,\xnz.mem_r_464_sv2v_reg ,\xnz.mem_r_463_sv2v_reg ,
  \xnz.mem_r_462_sv2v_reg ,\xnz.mem_r_461_sv2v_reg ,\xnz.mem_r_460_sv2v_reg ,
  \xnz.mem_r_459_sv2v_reg ,\xnz.mem_r_458_sv2v_reg ,\xnz.mem_r_457_sv2v_reg ,
  \xnz.mem_r_456_sv2v_reg ,\xnz.mem_r_455_sv2v_reg ,\xnz.mem_r_454_sv2v_reg ,\xnz.mem_r_453_sv2v_reg ,
  \xnz.mem_r_452_sv2v_reg ,\xnz.mem_r_451_sv2v_reg ,\xnz.mem_r_450_sv2v_reg ,
  \xnz.mem_r_449_sv2v_reg ,\xnz.mem_r_448_sv2v_reg ,\xnz.mem_r_447_sv2v_reg ,
  \xnz.mem_r_446_sv2v_reg ,\xnz.mem_r_445_sv2v_reg ,\xnz.mem_r_444_sv2v_reg ,
  \xnz.mem_r_443_sv2v_reg ,\xnz.mem_r_442_sv2v_reg ,\xnz.mem_r_441_sv2v_reg ,
  \xnz.mem_r_440_sv2v_reg ,\xnz.mem_r_439_sv2v_reg ,\xnz.mem_r_438_sv2v_reg ,\xnz.mem_r_437_sv2v_reg ,
  \xnz.mem_r_436_sv2v_reg ,\xnz.mem_r_435_sv2v_reg ,\xnz.mem_r_434_sv2v_reg ,
  \xnz.mem_r_433_sv2v_reg ,\xnz.mem_r_432_sv2v_reg ,\xnz.mem_r_431_sv2v_reg ,
  \xnz.mem_r_430_sv2v_reg ,\xnz.mem_r_429_sv2v_reg ,\xnz.mem_r_428_sv2v_reg ,
  \xnz.mem_r_427_sv2v_reg ,\xnz.mem_r_426_sv2v_reg ,\xnz.mem_r_425_sv2v_reg ,
  \xnz.mem_r_424_sv2v_reg ,\xnz.mem_r_423_sv2v_reg ,\xnz.mem_r_422_sv2v_reg ,\xnz.mem_r_421_sv2v_reg ,
  \xnz.mem_r_420_sv2v_reg ,\xnz.mem_r_419_sv2v_reg ,\xnz.mem_r_418_sv2v_reg ,
  \xnz.mem_r_417_sv2v_reg ,\xnz.mem_r_416_sv2v_reg ,\xnz.mem_r_415_sv2v_reg ,
  \xnz.mem_r_414_sv2v_reg ,\xnz.mem_r_413_sv2v_reg ,\xnz.mem_r_412_sv2v_reg ,
  \xnz.mem_r_411_sv2v_reg ,\xnz.mem_r_410_sv2v_reg ,\xnz.mem_r_409_sv2v_reg ,
  \xnz.mem_r_408_sv2v_reg ,\xnz.mem_r_407_sv2v_reg ,\xnz.mem_r_406_sv2v_reg ,\xnz.mem_r_405_sv2v_reg ,
  \xnz.mem_r_404_sv2v_reg ,\xnz.mem_r_403_sv2v_reg ,\xnz.mem_r_402_sv2v_reg ,
  \xnz.mem_r_401_sv2v_reg ,\xnz.mem_r_400_sv2v_reg ,\xnz.mem_r_399_sv2v_reg ,
  \xnz.mem_r_398_sv2v_reg ,\xnz.mem_r_397_sv2v_reg ,\xnz.mem_r_396_sv2v_reg ,
  \xnz.mem_r_395_sv2v_reg ,\xnz.mem_r_394_sv2v_reg ,\xnz.mem_r_393_sv2v_reg ,
  \xnz.mem_r_392_sv2v_reg ,\xnz.mem_r_391_sv2v_reg ,\xnz.mem_r_390_sv2v_reg ,\xnz.mem_r_389_sv2v_reg ,
  \xnz.mem_r_388_sv2v_reg ,\xnz.mem_r_387_sv2v_reg ,\xnz.mem_r_386_sv2v_reg ,
  \xnz.mem_r_385_sv2v_reg ,\xnz.mem_r_384_sv2v_reg ,\xnz.mem_r_383_sv2v_reg ,
  \xnz.mem_r_382_sv2v_reg ,\xnz.mem_r_381_sv2v_reg ,\xnz.mem_r_380_sv2v_reg ,
  \xnz.mem_r_379_sv2v_reg ,\xnz.mem_r_378_sv2v_reg ,\xnz.mem_r_377_sv2v_reg ,
  \xnz.mem_r_376_sv2v_reg ,\xnz.mem_r_375_sv2v_reg ,\xnz.mem_r_374_sv2v_reg ,\xnz.mem_r_373_sv2v_reg ,
  \xnz.mem_r_372_sv2v_reg ,\xnz.mem_r_371_sv2v_reg ,\xnz.mem_r_370_sv2v_reg ,
  \xnz.mem_r_369_sv2v_reg ,\xnz.mem_r_368_sv2v_reg ,\xnz.mem_r_367_sv2v_reg ,
  \xnz.mem_r_366_sv2v_reg ,\xnz.mem_r_365_sv2v_reg ,\xnz.mem_r_364_sv2v_reg ,
  \xnz.mem_r_363_sv2v_reg ,\xnz.mem_r_362_sv2v_reg ,\xnz.mem_r_361_sv2v_reg ,
  \xnz.mem_r_360_sv2v_reg ,\xnz.mem_r_359_sv2v_reg ,\xnz.mem_r_358_sv2v_reg ,\xnz.mem_r_357_sv2v_reg ,
  \xnz.mem_r_356_sv2v_reg ,\xnz.mem_r_355_sv2v_reg ,\xnz.mem_r_354_sv2v_reg ,
  \xnz.mem_r_353_sv2v_reg ,\xnz.mem_r_352_sv2v_reg ,\xnz.mem_r_351_sv2v_reg ,
  \xnz.mem_r_350_sv2v_reg ,\xnz.mem_r_349_sv2v_reg ,\xnz.mem_r_348_sv2v_reg ,
  \xnz.mem_r_347_sv2v_reg ,\xnz.mem_r_346_sv2v_reg ,\xnz.mem_r_345_sv2v_reg ,
  \xnz.mem_r_344_sv2v_reg ,\xnz.mem_r_343_sv2v_reg ,\xnz.mem_r_342_sv2v_reg ,\xnz.mem_r_341_sv2v_reg ,
  \xnz.mem_r_340_sv2v_reg ,\xnz.mem_r_339_sv2v_reg ,\xnz.mem_r_338_sv2v_reg ,
  \xnz.mem_r_337_sv2v_reg ,\xnz.mem_r_336_sv2v_reg ,\xnz.mem_r_335_sv2v_reg ,
  \xnz.mem_r_334_sv2v_reg ,\xnz.mem_r_333_sv2v_reg ,\xnz.mem_r_332_sv2v_reg ,
  \xnz.mem_r_331_sv2v_reg ,\xnz.mem_r_330_sv2v_reg ,\xnz.mem_r_329_sv2v_reg ,
  \xnz.mem_r_328_sv2v_reg ,\xnz.mem_r_327_sv2v_reg ,\xnz.mem_r_326_sv2v_reg ,\xnz.mem_r_325_sv2v_reg ,
  \xnz.mem_r_324_sv2v_reg ,\xnz.mem_r_323_sv2v_reg ,\xnz.mem_r_322_sv2v_reg ,
  \xnz.mem_r_321_sv2v_reg ,\xnz.mem_r_320_sv2v_reg ,\xnz.mem_r_319_sv2v_reg ,
  \xnz.mem_r_318_sv2v_reg ,\xnz.mem_r_317_sv2v_reg ,\xnz.mem_r_316_sv2v_reg ,
  \xnz.mem_r_315_sv2v_reg ,\xnz.mem_r_314_sv2v_reg ,\xnz.mem_r_313_sv2v_reg ,
  \xnz.mem_r_312_sv2v_reg ,\xnz.mem_r_311_sv2v_reg ,\xnz.mem_r_310_sv2v_reg ,\xnz.mem_r_309_sv2v_reg ,
  \xnz.mem_r_308_sv2v_reg ,\xnz.mem_r_307_sv2v_reg ,\xnz.mem_r_306_sv2v_reg ,
  \xnz.mem_r_305_sv2v_reg ,\xnz.mem_r_304_sv2v_reg ,\xnz.mem_r_303_sv2v_reg ,
  \xnz.mem_r_302_sv2v_reg ,\xnz.mem_r_301_sv2v_reg ,\xnz.mem_r_300_sv2v_reg ,
  \xnz.mem_r_299_sv2v_reg ,\xnz.mem_r_298_sv2v_reg ,\xnz.mem_r_297_sv2v_reg ,
  \xnz.mem_r_296_sv2v_reg ,\xnz.mem_r_295_sv2v_reg ,\xnz.mem_r_294_sv2v_reg ,\xnz.mem_r_293_sv2v_reg ,
  \xnz.mem_r_292_sv2v_reg ,\xnz.mem_r_291_sv2v_reg ,\xnz.mem_r_290_sv2v_reg ,
  \xnz.mem_r_289_sv2v_reg ,\xnz.mem_r_288_sv2v_reg ,\xnz.mem_r_287_sv2v_reg ,
  \xnz.mem_r_286_sv2v_reg ,\xnz.mem_r_285_sv2v_reg ,\xnz.mem_r_284_sv2v_reg ,
  \xnz.mem_r_283_sv2v_reg ,\xnz.mem_r_282_sv2v_reg ,\xnz.mem_r_281_sv2v_reg ,
  \xnz.mem_r_280_sv2v_reg ,\xnz.mem_r_279_sv2v_reg ,\xnz.mem_r_278_sv2v_reg ,\xnz.mem_r_277_sv2v_reg ,
  \xnz.mem_r_276_sv2v_reg ,\xnz.mem_r_275_sv2v_reg ,\xnz.mem_r_274_sv2v_reg ,
  \xnz.mem_r_273_sv2v_reg ,\xnz.mem_r_272_sv2v_reg ,\xnz.mem_r_271_sv2v_reg ,
  \xnz.mem_r_270_sv2v_reg ,\xnz.mem_r_269_sv2v_reg ,\xnz.mem_r_268_sv2v_reg ,
  \xnz.mem_r_267_sv2v_reg ,\xnz.mem_r_266_sv2v_reg ,\xnz.mem_r_265_sv2v_reg ,
  \xnz.mem_r_264_sv2v_reg ,\xnz.mem_r_263_sv2v_reg ,\xnz.mem_r_262_sv2v_reg ,\xnz.mem_r_261_sv2v_reg ,
  \xnz.mem_r_260_sv2v_reg ,\xnz.mem_r_259_sv2v_reg ,\xnz.mem_r_258_sv2v_reg ,
  \xnz.mem_r_257_sv2v_reg ,\xnz.mem_r_256_sv2v_reg ,\xnz.mem_r_255_sv2v_reg ,
  \xnz.mem_r_254_sv2v_reg ,\xnz.mem_r_253_sv2v_reg ,\xnz.mem_r_252_sv2v_reg ,
  \xnz.mem_r_251_sv2v_reg ,\xnz.mem_r_250_sv2v_reg ,\xnz.mem_r_249_sv2v_reg ,
  \xnz.mem_r_248_sv2v_reg ,\xnz.mem_r_247_sv2v_reg ,\xnz.mem_r_246_sv2v_reg ,\xnz.mem_r_245_sv2v_reg ,
  \xnz.mem_r_244_sv2v_reg ,\xnz.mem_r_243_sv2v_reg ,\xnz.mem_r_242_sv2v_reg ,
  \xnz.mem_r_241_sv2v_reg ,\xnz.mem_r_240_sv2v_reg ,\xnz.mem_r_239_sv2v_reg ,
  \xnz.mem_r_238_sv2v_reg ,\xnz.mem_r_237_sv2v_reg ,\xnz.mem_r_236_sv2v_reg ,
  \xnz.mem_r_235_sv2v_reg ,\xnz.mem_r_234_sv2v_reg ,\xnz.mem_r_233_sv2v_reg ,
  \xnz.mem_r_232_sv2v_reg ,\xnz.mem_r_231_sv2v_reg ,\xnz.mem_r_230_sv2v_reg ,\xnz.mem_r_229_sv2v_reg ,
  \xnz.mem_r_228_sv2v_reg ,\xnz.mem_r_227_sv2v_reg ,\xnz.mem_r_226_sv2v_reg ,
  \xnz.mem_r_225_sv2v_reg ,\xnz.mem_r_224_sv2v_reg ,\xnz.mem_r_223_sv2v_reg ,
  \xnz.mem_r_222_sv2v_reg ,\xnz.mem_r_221_sv2v_reg ,\xnz.mem_r_220_sv2v_reg ,
  \xnz.mem_r_219_sv2v_reg ,\xnz.mem_r_218_sv2v_reg ,\xnz.mem_r_217_sv2v_reg ,
  \xnz.mem_r_216_sv2v_reg ,\xnz.mem_r_215_sv2v_reg ,\xnz.mem_r_214_sv2v_reg ,\xnz.mem_r_213_sv2v_reg ,
  \xnz.mem_r_212_sv2v_reg ,\xnz.mem_r_211_sv2v_reg ,\xnz.mem_r_210_sv2v_reg ,
  \xnz.mem_r_209_sv2v_reg ,\xnz.mem_r_208_sv2v_reg ,\xnz.mem_r_207_sv2v_reg ,
  \xnz.mem_r_206_sv2v_reg ,\xnz.mem_r_205_sv2v_reg ,\xnz.mem_r_204_sv2v_reg ,
  \xnz.mem_r_203_sv2v_reg ,\xnz.mem_r_202_sv2v_reg ,\xnz.mem_r_201_sv2v_reg ,
  \xnz.mem_r_200_sv2v_reg ,\xnz.mem_r_199_sv2v_reg ,\xnz.mem_r_198_sv2v_reg ,\xnz.mem_r_197_sv2v_reg ,
  \xnz.mem_r_196_sv2v_reg ,\xnz.mem_r_195_sv2v_reg ,\xnz.mem_r_194_sv2v_reg ,
  \xnz.mem_r_193_sv2v_reg ,\xnz.mem_r_192_sv2v_reg ,\xnz.mem_r_191_sv2v_reg ,
  \xnz.mem_r_190_sv2v_reg ,\xnz.mem_r_189_sv2v_reg ,\xnz.mem_r_188_sv2v_reg ,
  \xnz.mem_r_187_sv2v_reg ,\xnz.mem_r_186_sv2v_reg ,\xnz.mem_r_185_sv2v_reg ,
  \xnz.mem_r_184_sv2v_reg ,\xnz.mem_r_183_sv2v_reg ,\xnz.mem_r_182_sv2v_reg ,\xnz.mem_r_181_sv2v_reg ,
  \xnz.mem_r_180_sv2v_reg ,\xnz.mem_r_179_sv2v_reg ,\xnz.mem_r_178_sv2v_reg ,
  \xnz.mem_r_177_sv2v_reg ,\xnz.mem_r_176_sv2v_reg ,\xnz.mem_r_175_sv2v_reg ,
  \xnz.mem_r_174_sv2v_reg ,\xnz.mem_r_173_sv2v_reg ,\xnz.mem_r_172_sv2v_reg ,
  \xnz.mem_r_171_sv2v_reg ,\xnz.mem_r_170_sv2v_reg ,\xnz.mem_r_169_sv2v_reg ,
  \xnz.mem_r_168_sv2v_reg ,\xnz.mem_r_167_sv2v_reg ,\xnz.mem_r_166_sv2v_reg ,\xnz.mem_r_165_sv2v_reg ,
  \xnz.mem_r_164_sv2v_reg ,\xnz.mem_r_163_sv2v_reg ,\xnz.mem_r_162_sv2v_reg ,
  \xnz.mem_r_161_sv2v_reg ,\xnz.mem_r_160_sv2v_reg ,\xnz.mem_r_159_sv2v_reg ,
  \xnz.mem_r_158_sv2v_reg ,\xnz.mem_r_157_sv2v_reg ,\xnz.mem_r_156_sv2v_reg ,
  \xnz.mem_r_155_sv2v_reg ,\xnz.mem_r_154_sv2v_reg ,\xnz.mem_r_153_sv2v_reg ,
  \xnz.mem_r_152_sv2v_reg ,\xnz.mem_r_151_sv2v_reg ,\xnz.mem_r_150_sv2v_reg ,\xnz.mem_r_149_sv2v_reg ,
  \xnz.mem_r_148_sv2v_reg ,\xnz.mem_r_147_sv2v_reg ,\xnz.mem_r_146_sv2v_reg ,
  \xnz.mem_r_145_sv2v_reg ,\xnz.mem_r_144_sv2v_reg ,\xnz.mem_r_143_sv2v_reg ,
  \xnz.mem_r_142_sv2v_reg ,\xnz.mem_r_141_sv2v_reg ,\xnz.mem_r_140_sv2v_reg ,
  \xnz.mem_r_139_sv2v_reg ,\xnz.mem_r_138_sv2v_reg ,\xnz.mem_r_137_sv2v_reg ,
  \xnz.mem_r_136_sv2v_reg ,\xnz.mem_r_135_sv2v_reg ,\xnz.mem_r_134_sv2v_reg ,\xnz.mem_r_133_sv2v_reg ,
  \xnz.mem_r_132_sv2v_reg ,\xnz.mem_r_131_sv2v_reg ,\xnz.mem_r_130_sv2v_reg ,
  \xnz.mem_r_129_sv2v_reg ,\xnz.mem_r_128_sv2v_reg ,\xnz.mem_r_127_sv2v_reg ,
  \xnz.mem_r_126_sv2v_reg ,\xnz.mem_r_125_sv2v_reg ,\xnz.mem_r_124_sv2v_reg ,
  \xnz.mem_r_123_sv2v_reg ,\xnz.mem_r_122_sv2v_reg ,\xnz.mem_r_121_sv2v_reg ,
  \xnz.mem_r_120_sv2v_reg ,\xnz.mem_r_119_sv2v_reg ,\xnz.mem_r_118_sv2v_reg ,\xnz.mem_r_117_sv2v_reg ,
  \xnz.mem_r_116_sv2v_reg ,\xnz.mem_r_115_sv2v_reg ,\xnz.mem_r_114_sv2v_reg ,
  \xnz.mem_r_113_sv2v_reg ,\xnz.mem_r_112_sv2v_reg ,\xnz.mem_r_111_sv2v_reg ,
  \xnz.mem_r_110_sv2v_reg ,\xnz.mem_r_109_sv2v_reg ,\xnz.mem_r_108_sv2v_reg ,
  \xnz.mem_r_107_sv2v_reg ,\xnz.mem_r_106_sv2v_reg ,\xnz.mem_r_105_sv2v_reg ,
  \xnz.mem_r_104_sv2v_reg ,\xnz.mem_r_103_sv2v_reg ,\xnz.mem_r_102_sv2v_reg ,\xnz.mem_r_101_sv2v_reg ,
  \xnz.mem_r_100_sv2v_reg ,\xnz.mem_r_99_sv2v_reg ,\xnz.mem_r_98_sv2v_reg ,
  \xnz.mem_r_97_sv2v_reg ,\xnz.mem_r_96_sv2v_reg ,\xnz.mem_r_95_sv2v_reg ,
  \xnz.mem_r_94_sv2v_reg ,\xnz.mem_r_93_sv2v_reg ,\xnz.mem_r_92_sv2v_reg ,\xnz.mem_r_91_sv2v_reg ,
  \xnz.mem_r_90_sv2v_reg ,\xnz.mem_r_89_sv2v_reg ,\xnz.mem_r_88_sv2v_reg ,
  \xnz.mem_r_87_sv2v_reg ,\xnz.mem_r_86_sv2v_reg ,\xnz.mem_r_85_sv2v_reg ,
  \xnz.mem_r_84_sv2v_reg ,\xnz.mem_r_83_sv2v_reg ,\xnz.mem_r_82_sv2v_reg ,\xnz.mem_r_81_sv2v_reg ,
  \xnz.mem_r_80_sv2v_reg ,\xnz.mem_r_79_sv2v_reg ,\xnz.mem_r_78_sv2v_reg ,
  \xnz.mem_r_77_sv2v_reg ,\xnz.mem_r_76_sv2v_reg ,\xnz.mem_r_75_sv2v_reg ,
  \xnz.mem_r_74_sv2v_reg ,\xnz.mem_r_73_sv2v_reg ,\xnz.mem_r_72_sv2v_reg ,\xnz.mem_r_71_sv2v_reg ,
  \xnz.mem_r_70_sv2v_reg ,\xnz.mem_r_69_sv2v_reg ,\xnz.mem_r_68_sv2v_reg ,
  \xnz.mem_r_67_sv2v_reg ,\xnz.mem_r_66_sv2v_reg ,\xnz.mem_r_65_sv2v_reg ,
  \xnz.mem_r_64_sv2v_reg ,\xnz.mem_r_63_sv2v_reg ,\xnz.mem_r_62_sv2v_reg ,\xnz.mem_r_61_sv2v_reg ,
  \xnz.mem_r_60_sv2v_reg ,\xnz.mem_r_59_sv2v_reg ,\xnz.mem_r_58_sv2v_reg ,
  \xnz.mem_r_57_sv2v_reg ,\xnz.mem_r_56_sv2v_reg ,\xnz.mem_r_55_sv2v_reg ,
  \xnz.mem_r_54_sv2v_reg ,\xnz.mem_r_53_sv2v_reg ,\xnz.mem_r_52_sv2v_reg ,\xnz.mem_r_51_sv2v_reg ,
  \xnz.mem_r_50_sv2v_reg ,\xnz.mem_r_49_sv2v_reg ,\xnz.mem_r_48_sv2v_reg ,
  \xnz.mem_r_47_sv2v_reg ,\xnz.mem_r_46_sv2v_reg ,\xnz.mem_r_45_sv2v_reg ,
  \xnz.mem_r_44_sv2v_reg ,\xnz.mem_r_43_sv2v_reg ,\xnz.mem_r_42_sv2v_reg ,\xnz.mem_r_41_sv2v_reg ,
  \xnz.mem_r_40_sv2v_reg ,\xnz.mem_r_39_sv2v_reg ,\xnz.mem_r_38_sv2v_reg ,
  \xnz.mem_r_37_sv2v_reg ,\xnz.mem_r_36_sv2v_reg ,\xnz.mem_r_35_sv2v_reg ,
  \xnz.mem_r_34_sv2v_reg ,\xnz.mem_r_33_sv2v_reg ,\xnz.mem_r_32_sv2v_reg ,\xnz.mem_r_31_sv2v_reg ,
  \xnz.mem_r_30_sv2v_reg ,\xnz.mem_r_29_sv2v_reg ,\xnz.mem_r_28_sv2v_reg ,
  \xnz.mem_r_27_sv2v_reg ,\xnz.mem_r_26_sv2v_reg ,\xnz.mem_r_25_sv2v_reg ,
  \xnz.mem_r_24_sv2v_reg ,\xnz.mem_r_23_sv2v_reg ,\xnz.mem_r_22_sv2v_reg ,\xnz.mem_r_21_sv2v_reg ,
  \xnz.mem_r_20_sv2v_reg ,\xnz.mem_r_19_sv2v_reg ,\xnz.mem_r_18_sv2v_reg ,
  \xnz.mem_r_17_sv2v_reg ,\xnz.mem_r_16_sv2v_reg ,\xnz.mem_r_15_sv2v_reg ,
  \xnz.mem_r_14_sv2v_reg ,\xnz.mem_r_13_sv2v_reg ,\xnz.mem_r_12_sv2v_reg ,\xnz.mem_r_11_sv2v_reg ,
  \xnz.mem_r_10_sv2v_reg ,\xnz.mem_r_9_sv2v_reg ,\xnz.mem_r_8_sv2v_reg ,
  \xnz.mem_r_7_sv2v_reg ,\xnz.mem_r_6_sv2v_reg ,\xnz.mem_r_5_sv2v_reg ,\xnz.mem_r_4_sv2v_reg ,
  \xnz.mem_r_3_sv2v_reg ,\xnz.mem_r_2_sv2v_reg ,\xnz.mem_r_1_sv2v_reg ,
  \xnz.mem_r_0_sv2v_reg ;
  assign r_addr_r[14] = r_addr_r_14_sv2v_reg;
  assign r_addr_r[13] = r_addr_r_13_sv2v_reg;
  assign r_addr_r[12] = r_addr_r_12_sv2v_reg;
  assign r_addr_r[11] = r_addr_r_11_sv2v_reg;
  assign r_addr_r[10] = r_addr_r_10_sv2v_reg;
  assign r_addr_r[9] = r_addr_r_9_sv2v_reg;
  assign r_addr_r[8] = r_addr_r_8_sv2v_reg;
  assign r_addr_r[7] = r_addr_r_7_sv2v_reg;
  assign r_addr_r[6] = r_addr_r_6_sv2v_reg;
  assign r_addr_r[5] = r_addr_r_5_sv2v_reg;
  assign r_addr_r[4] = r_addr_r_4_sv2v_reg;
  assign r_addr_r[3] = r_addr_r_3_sv2v_reg;
  assign r_addr_r[2] = r_addr_r_2_sv2v_reg;
  assign r_addr_r[1] = r_addr_r_1_sv2v_reg;
  assign r_addr_r[0] = r_addr_r_0_sv2v_reg;
  assign \xnz.mem_r [1055] = \xnz.mem_r_1055_sv2v_reg ;
  assign \xnz.mem_r [1054] = \xnz.mem_r_1054_sv2v_reg ;
  assign \xnz.mem_r [1053] = \xnz.mem_r_1053_sv2v_reg ;
  assign \xnz.mem_r [1052] = \xnz.mem_r_1052_sv2v_reg ;
  assign \xnz.mem_r [1051] = \xnz.mem_r_1051_sv2v_reg ;
  assign \xnz.mem_r [1050] = \xnz.mem_r_1050_sv2v_reg ;
  assign \xnz.mem_r [1049] = \xnz.mem_r_1049_sv2v_reg ;
  assign \xnz.mem_r [1048] = \xnz.mem_r_1048_sv2v_reg ;
  assign \xnz.mem_r [1047] = \xnz.mem_r_1047_sv2v_reg ;
  assign \xnz.mem_r [1046] = \xnz.mem_r_1046_sv2v_reg ;
  assign \xnz.mem_r [1045] = \xnz.mem_r_1045_sv2v_reg ;
  assign \xnz.mem_r [1044] = \xnz.mem_r_1044_sv2v_reg ;
  assign \xnz.mem_r [1043] = \xnz.mem_r_1043_sv2v_reg ;
  assign \xnz.mem_r [1042] = \xnz.mem_r_1042_sv2v_reg ;
  assign \xnz.mem_r [1041] = \xnz.mem_r_1041_sv2v_reg ;
  assign \xnz.mem_r [1040] = \xnz.mem_r_1040_sv2v_reg ;
  assign \xnz.mem_r [1039] = \xnz.mem_r_1039_sv2v_reg ;
  assign \xnz.mem_r [1038] = \xnz.mem_r_1038_sv2v_reg ;
  assign \xnz.mem_r [1037] = \xnz.mem_r_1037_sv2v_reg ;
  assign \xnz.mem_r [1036] = \xnz.mem_r_1036_sv2v_reg ;
  assign \xnz.mem_r [1035] = \xnz.mem_r_1035_sv2v_reg ;
  assign \xnz.mem_r [1034] = \xnz.mem_r_1034_sv2v_reg ;
  assign \xnz.mem_r [1033] = \xnz.mem_r_1033_sv2v_reg ;
  assign \xnz.mem_r [1032] = \xnz.mem_r_1032_sv2v_reg ;
  assign \xnz.mem_r [1031] = \xnz.mem_r_1031_sv2v_reg ;
  assign \xnz.mem_r [1030] = \xnz.mem_r_1030_sv2v_reg ;
  assign \xnz.mem_r [1029] = \xnz.mem_r_1029_sv2v_reg ;
  assign \xnz.mem_r [1028] = \xnz.mem_r_1028_sv2v_reg ;
  assign \xnz.mem_r [1027] = \xnz.mem_r_1027_sv2v_reg ;
  assign \xnz.mem_r [1026] = \xnz.mem_r_1026_sv2v_reg ;
  assign \xnz.mem_r [1025] = \xnz.mem_r_1025_sv2v_reg ;
  assign \xnz.mem_r [1024] = \xnz.mem_r_1024_sv2v_reg ;
  assign \xnz.mem_r [1023] = \xnz.mem_r_1023_sv2v_reg ;
  assign \xnz.mem_r [1022] = \xnz.mem_r_1022_sv2v_reg ;
  assign \xnz.mem_r [1021] = \xnz.mem_r_1021_sv2v_reg ;
  assign \xnz.mem_r [1020] = \xnz.mem_r_1020_sv2v_reg ;
  assign \xnz.mem_r [1019] = \xnz.mem_r_1019_sv2v_reg ;
  assign \xnz.mem_r [1018] = \xnz.mem_r_1018_sv2v_reg ;
  assign \xnz.mem_r [1017] = \xnz.mem_r_1017_sv2v_reg ;
  assign \xnz.mem_r [1016] = \xnz.mem_r_1016_sv2v_reg ;
  assign \xnz.mem_r [1015] = \xnz.mem_r_1015_sv2v_reg ;
  assign \xnz.mem_r [1014] = \xnz.mem_r_1014_sv2v_reg ;
  assign \xnz.mem_r [1013] = \xnz.mem_r_1013_sv2v_reg ;
  assign \xnz.mem_r [1012] = \xnz.mem_r_1012_sv2v_reg ;
  assign \xnz.mem_r [1011] = \xnz.mem_r_1011_sv2v_reg ;
  assign \xnz.mem_r [1010] = \xnz.mem_r_1010_sv2v_reg ;
  assign \xnz.mem_r [1009] = \xnz.mem_r_1009_sv2v_reg ;
  assign \xnz.mem_r [1008] = \xnz.mem_r_1008_sv2v_reg ;
  assign \xnz.mem_r [1007] = \xnz.mem_r_1007_sv2v_reg ;
  assign \xnz.mem_r [1006] = \xnz.mem_r_1006_sv2v_reg ;
  assign \xnz.mem_r [1005] = \xnz.mem_r_1005_sv2v_reg ;
  assign \xnz.mem_r [1004] = \xnz.mem_r_1004_sv2v_reg ;
  assign \xnz.mem_r [1003] = \xnz.mem_r_1003_sv2v_reg ;
  assign \xnz.mem_r [1002] = \xnz.mem_r_1002_sv2v_reg ;
  assign \xnz.mem_r [1001] = \xnz.mem_r_1001_sv2v_reg ;
  assign \xnz.mem_r [1000] = \xnz.mem_r_1000_sv2v_reg ;
  assign \xnz.mem_r [999] = \xnz.mem_r_999_sv2v_reg ;
  assign \xnz.mem_r [998] = \xnz.mem_r_998_sv2v_reg ;
  assign \xnz.mem_r [997] = \xnz.mem_r_997_sv2v_reg ;
  assign \xnz.mem_r [996] = \xnz.mem_r_996_sv2v_reg ;
  assign \xnz.mem_r [995] = \xnz.mem_r_995_sv2v_reg ;
  assign \xnz.mem_r [994] = \xnz.mem_r_994_sv2v_reg ;
  assign \xnz.mem_r [993] = \xnz.mem_r_993_sv2v_reg ;
  assign \xnz.mem_r [992] = \xnz.mem_r_992_sv2v_reg ;
  assign \xnz.mem_r [991] = \xnz.mem_r_991_sv2v_reg ;
  assign \xnz.mem_r [990] = \xnz.mem_r_990_sv2v_reg ;
  assign \xnz.mem_r [989] = \xnz.mem_r_989_sv2v_reg ;
  assign \xnz.mem_r [988] = \xnz.mem_r_988_sv2v_reg ;
  assign \xnz.mem_r [987] = \xnz.mem_r_987_sv2v_reg ;
  assign \xnz.mem_r [986] = \xnz.mem_r_986_sv2v_reg ;
  assign \xnz.mem_r [985] = \xnz.mem_r_985_sv2v_reg ;
  assign \xnz.mem_r [984] = \xnz.mem_r_984_sv2v_reg ;
  assign \xnz.mem_r [983] = \xnz.mem_r_983_sv2v_reg ;
  assign \xnz.mem_r [982] = \xnz.mem_r_982_sv2v_reg ;
  assign \xnz.mem_r [981] = \xnz.mem_r_981_sv2v_reg ;
  assign \xnz.mem_r [980] = \xnz.mem_r_980_sv2v_reg ;
  assign \xnz.mem_r [979] = \xnz.mem_r_979_sv2v_reg ;
  assign \xnz.mem_r [978] = \xnz.mem_r_978_sv2v_reg ;
  assign \xnz.mem_r [977] = \xnz.mem_r_977_sv2v_reg ;
  assign \xnz.mem_r [976] = \xnz.mem_r_976_sv2v_reg ;
  assign \xnz.mem_r [975] = \xnz.mem_r_975_sv2v_reg ;
  assign \xnz.mem_r [974] = \xnz.mem_r_974_sv2v_reg ;
  assign \xnz.mem_r [973] = \xnz.mem_r_973_sv2v_reg ;
  assign \xnz.mem_r [972] = \xnz.mem_r_972_sv2v_reg ;
  assign \xnz.mem_r [971] = \xnz.mem_r_971_sv2v_reg ;
  assign \xnz.mem_r [970] = \xnz.mem_r_970_sv2v_reg ;
  assign \xnz.mem_r [969] = \xnz.mem_r_969_sv2v_reg ;
  assign \xnz.mem_r [968] = \xnz.mem_r_968_sv2v_reg ;
  assign \xnz.mem_r [967] = \xnz.mem_r_967_sv2v_reg ;
  assign \xnz.mem_r [966] = \xnz.mem_r_966_sv2v_reg ;
  assign \xnz.mem_r [965] = \xnz.mem_r_965_sv2v_reg ;
  assign \xnz.mem_r [964] = \xnz.mem_r_964_sv2v_reg ;
  assign \xnz.mem_r [963] = \xnz.mem_r_963_sv2v_reg ;
  assign \xnz.mem_r [962] = \xnz.mem_r_962_sv2v_reg ;
  assign \xnz.mem_r [961] = \xnz.mem_r_961_sv2v_reg ;
  assign \xnz.mem_r [960] = \xnz.mem_r_960_sv2v_reg ;
  assign \xnz.mem_r [959] = \xnz.mem_r_959_sv2v_reg ;
  assign \xnz.mem_r [958] = \xnz.mem_r_958_sv2v_reg ;
  assign \xnz.mem_r [957] = \xnz.mem_r_957_sv2v_reg ;
  assign \xnz.mem_r [956] = \xnz.mem_r_956_sv2v_reg ;
  assign \xnz.mem_r [955] = \xnz.mem_r_955_sv2v_reg ;
  assign \xnz.mem_r [954] = \xnz.mem_r_954_sv2v_reg ;
  assign \xnz.mem_r [953] = \xnz.mem_r_953_sv2v_reg ;
  assign \xnz.mem_r [952] = \xnz.mem_r_952_sv2v_reg ;
  assign \xnz.mem_r [951] = \xnz.mem_r_951_sv2v_reg ;
  assign \xnz.mem_r [950] = \xnz.mem_r_950_sv2v_reg ;
  assign \xnz.mem_r [949] = \xnz.mem_r_949_sv2v_reg ;
  assign \xnz.mem_r [948] = \xnz.mem_r_948_sv2v_reg ;
  assign \xnz.mem_r [947] = \xnz.mem_r_947_sv2v_reg ;
  assign \xnz.mem_r [946] = \xnz.mem_r_946_sv2v_reg ;
  assign \xnz.mem_r [945] = \xnz.mem_r_945_sv2v_reg ;
  assign \xnz.mem_r [944] = \xnz.mem_r_944_sv2v_reg ;
  assign \xnz.mem_r [943] = \xnz.mem_r_943_sv2v_reg ;
  assign \xnz.mem_r [942] = \xnz.mem_r_942_sv2v_reg ;
  assign \xnz.mem_r [941] = \xnz.mem_r_941_sv2v_reg ;
  assign \xnz.mem_r [940] = \xnz.mem_r_940_sv2v_reg ;
  assign \xnz.mem_r [939] = \xnz.mem_r_939_sv2v_reg ;
  assign \xnz.mem_r [938] = \xnz.mem_r_938_sv2v_reg ;
  assign \xnz.mem_r [937] = \xnz.mem_r_937_sv2v_reg ;
  assign \xnz.mem_r [936] = \xnz.mem_r_936_sv2v_reg ;
  assign \xnz.mem_r [935] = \xnz.mem_r_935_sv2v_reg ;
  assign \xnz.mem_r [934] = \xnz.mem_r_934_sv2v_reg ;
  assign \xnz.mem_r [933] = \xnz.mem_r_933_sv2v_reg ;
  assign \xnz.mem_r [932] = \xnz.mem_r_932_sv2v_reg ;
  assign \xnz.mem_r [931] = \xnz.mem_r_931_sv2v_reg ;
  assign \xnz.mem_r [930] = \xnz.mem_r_930_sv2v_reg ;
  assign \xnz.mem_r [929] = \xnz.mem_r_929_sv2v_reg ;
  assign \xnz.mem_r [928] = \xnz.mem_r_928_sv2v_reg ;
  assign \xnz.mem_r [927] = \xnz.mem_r_927_sv2v_reg ;
  assign \xnz.mem_r [926] = \xnz.mem_r_926_sv2v_reg ;
  assign \xnz.mem_r [925] = \xnz.mem_r_925_sv2v_reg ;
  assign \xnz.mem_r [924] = \xnz.mem_r_924_sv2v_reg ;
  assign \xnz.mem_r [923] = \xnz.mem_r_923_sv2v_reg ;
  assign \xnz.mem_r [922] = \xnz.mem_r_922_sv2v_reg ;
  assign \xnz.mem_r [921] = \xnz.mem_r_921_sv2v_reg ;
  assign \xnz.mem_r [920] = \xnz.mem_r_920_sv2v_reg ;
  assign \xnz.mem_r [919] = \xnz.mem_r_919_sv2v_reg ;
  assign \xnz.mem_r [918] = \xnz.mem_r_918_sv2v_reg ;
  assign \xnz.mem_r [917] = \xnz.mem_r_917_sv2v_reg ;
  assign \xnz.mem_r [916] = \xnz.mem_r_916_sv2v_reg ;
  assign \xnz.mem_r [915] = \xnz.mem_r_915_sv2v_reg ;
  assign \xnz.mem_r [914] = \xnz.mem_r_914_sv2v_reg ;
  assign \xnz.mem_r [913] = \xnz.mem_r_913_sv2v_reg ;
  assign \xnz.mem_r [912] = \xnz.mem_r_912_sv2v_reg ;
  assign \xnz.mem_r [911] = \xnz.mem_r_911_sv2v_reg ;
  assign \xnz.mem_r [910] = \xnz.mem_r_910_sv2v_reg ;
  assign \xnz.mem_r [909] = \xnz.mem_r_909_sv2v_reg ;
  assign \xnz.mem_r [908] = \xnz.mem_r_908_sv2v_reg ;
  assign \xnz.mem_r [907] = \xnz.mem_r_907_sv2v_reg ;
  assign \xnz.mem_r [906] = \xnz.mem_r_906_sv2v_reg ;
  assign \xnz.mem_r [905] = \xnz.mem_r_905_sv2v_reg ;
  assign \xnz.mem_r [904] = \xnz.mem_r_904_sv2v_reg ;
  assign \xnz.mem_r [903] = \xnz.mem_r_903_sv2v_reg ;
  assign \xnz.mem_r [902] = \xnz.mem_r_902_sv2v_reg ;
  assign \xnz.mem_r [901] = \xnz.mem_r_901_sv2v_reg ;
  assign \xnz.mem_r [900] = \xnz.mem_r_900_sv2v_reg ;
  assign \xnz.mem_r [899] = \xnz.mem_r_899_sv2v_reg ;
  assign \xnz.mem_r [898] = \xnz.mem_r_898_sv2v_reg ;
  assign \xnz.mem_r [897] = \xnz.mem_r_897_sv2v_reg ;
  assign \xnz.mem_r [896] = \xnz.mem_r_896_sv2v_reg ;
  assign \xnz.mem_r [895] = \xnz.mem_r_895_sv2v_reg ;
  assign \xnz.mem_r [894] = \xnz.mem_r_894_sv2v_reg ;
  assign \xnz.mem_r [893] = \xnz.mem_r_893_sv2v_reg ;
  assign \xnz.mem_r [892] = \xnz.mem_r_892_sv2v_reg ;
  assign \xnz.mem_r [891] = \xnz.mem_r_891_sv2v_reg ;
  assign \xnz.mem_r [890] = \xnz.mem_r_890_sv2v_reg ;
  assign \xnz.mem_r [889] = \xnz.mem_r_889_sv2v_reg ;
  assign \xnz.mem_r [888] = \xnz.mem_r_888_sv2v_reg ;
  assign \xnz.mem_r [887] = \xnz.mem_r_887_sv2v_reg ;
  assign \xnz.mem_r [886] = \xnz.mem_r_886_sv2v_reg ;
  assign \xnz.mem_r [885] = \xnz.mem_r_885_sv2v_reg ;
  assign \xnz.mem_r [884] = \xnz.mem_r_884_sv2v_reg ;
  assign \xnz.mem_r [883] = \xnz.mem_r_883_sv2v_reg ;
  assign \xnz.mem_r [882] = \xnz.mem_r_882_sv2v_reg ;
  assign \xnz.mem_r [881] = \xnz.mem_r_881_sv2v_reg ;
  assign \xnz.mem_r [880] = \xnz.mem_r_880_sv2v_reg ;
  assign \xnz.mem_r [879] = \xnz.mem_r_879_sv2v_reg ;
  assign \xnz.mem_r [878] = \xnz.mem_r_878_sv2v_reg ;
  assign \xnz.mem_r [877] = \xnz.mem_r_877_sv2v_reg ;
  assign \xnz.mem_r [876] = \xnz.mem_r_876_sv2v_reg ;
  assign \xnz.mem_r [875] = \xnz.mem_r_875_sv2v_reg ;
  assign \xnz.mem_r [874] = \xnz.mem_r_874_sv2v_reg ;
  assign \xnz.mem_r [873] = \xnz.mem_r_873_sv2v_reg ;
  assign \xnz.mem_r [872] = \xnz.mem_r_872_sv2v_reg ;
  assign \xnz.mem_r [871] = \xnz.mem_r_871_sv2v_reg ;
  assign \xnz.mem_r [870] = \xnz.mem_r_870_sv2v_reg ;
  assign \xnz.mem_r [869] = \xnz.mem_r_869_sv2v_reg ;
  assign \xnz.mem_r [868] = \xnz.mem_r_868_sv2v_reg ;
  assign \xnz.mem_r [867] = \xnz.mem_r_867_sv2v_reg ;
  assign \xnz.mem_r [866] = \xnz.mem_r_866_sv2v_reg ;
  assign \xnz.mem_r [865] = \xnz.mem_r_865_sv2v_reg ;
  assign \xnz.mem_r [864] = \xnz.mem_r_864_sv2v_reg ;
  assign \xnz.mem_r [863] = \xnz.mem_r_863_sv2v_reg ;
  assign \xnz.mem_r [862] = \xnz.mem_r_862_sv2v_reg ;
  assign \xnz.mem_r [861] = \xnz.mem_r_861_sv2v_reg ;
  assign \xnz.mem_r [860] = \xnz.mem_r_860_sv2v_reg ;
  assign \xnz.mem_r [859] = \xnz.mem_r_859_sv2v_reg ;
  assign \xnz.mem_r [858] = \xnz.mem_r_858_sv2v_reg ;
  assign \xnz.mem_r [857] = \xnz.mem_r_857_sv2v_reg ;
  assign \xnz.mem_r [856] = \xnz.mem_r_856_sv2v_reg ;
  assign \xnz.mem_r [855] = \xnz.mem_r_855_sv2v_reg ;
  assign \xnz.mem_r [854] = \xnz.mem_r_854_sv2v_reg ;
  assign \xnz.mem_r [853] = \xnz.mem_r_853_sv2v_reg ;
  assign \xnz.mem_r [852] = \xnz.mem_r_852_sv2v_reg ;
  assign \xnz.mem_r [851] = \xnz.mem_r_851_sv2v_reg ;
  assign \xnz.mem_r [850] = \xnz.mem_r_850_sv2v_reg ;
  assign \xnz.mem_r [849] = \xnz.mem_r_849_sv2v_reg ;
  assign \xnz.mem_r [848] = \xnz.mem_r_848_sv2v_reg ;
  assign \xnz.mem_r [847] = \xnz.mem_r_847_sv2v_reg ;
  assign \xnz.mem_r [846] = \xnz.mem_r_846_sv2v_reg ;
  assign \xnz.mem_r [845] = \xnz.mem_r_845_sv2v_reg ;
  assign \xnz.mem_r [844] = \xnz.mem_r_844_sv2v_reg ;
  assign \xnz.mem_r [843] = \xnz.mem_r_843_sv2v_reg ;
  assign \xnz.mem_r [842] = \xnz.mem_r_842_sv2v_reg ;
  assign \xnz.mem_r [841] = \xnz.mem_r_841_sv2v_reg ;
  assign \xnz.mem_r [840] = \xnz.mem_r_840_sv2v_reg ;
  assign \xnz.mem_r [839] = \xnz.mem_r_839_sv2v_reg ;
  assign \xnz.mem_r [838] = \xnz.mem_r_838_sv2v_reg ;
  assign \xnz.mem_r [837] = \xnz.mem_r_837_sv2v_reg ;
  assign \xnz.mem_r [836] = \xnz.mem_r_836_sv2v_reg ;
  assign \xnz.mem_r [835] = \xnz.mem_r_835_sv2v_reg ;
  assign \xnz.mem_r [834] = \xnz.mem_r_834_sv2v_reg ;
  assign \xnz.mem_r [833] = \xnz.mem_r_833_sv2v_reg ;
  assign \xnz.mem_r [832] = \xnz.mem_r_832_sv2v_reg ;
  assign \xnz.mem_r [831] = \xnz.mem_r_831_sv2v_reg ;
  assign \xnz.mem_r [830] = \xnz.mem_r_830_sv2v_reg ;
  assign \xnz.mem_r [829] = \xnz.mem_r_829_sv2v_reg ;
  assign \xnz.mem_r [828] = \xnz.mem_r_828_sv2v_reg ;
  assign \xnz.mem_r [827] = \xnz.mem_r_827_sv2v_reg ;
  assign \xnz.mem_r [826] = \xnz.mem_r_826_sv2v_reg ;
  assign \xnz.mem_r [825] = \xnz.mem_r_825_sv2v_reg ;
  assign \xnz.mem_r [824] = \xnz.mem_r_824_sv2v_reg ;
  assign \xnz.mem_r [823] = \xnz.mem_r_823_sv2v_reg ;
  assign \xnz.mem_r [822] = \xnz.mem_r_822_sv2v_reg ;
  assign \xnz.mem_r [821] = \xnz.mem_r_821_sv2v_reg ;
  assign \xnz.mem_r [820] = \xnz.mem_r_820_sv2v_reg ;
  assign \xnz.mem_r [819] = \xnz.mem_r_819_sv2v_reg ;
  assign \xnz.mem_r [818] = \xnz.mem_r_818_sv2v_reg ;
  assign \xnz.mem_r [817] = \xnz.mem_r_817_sv2v_reg ;
  assign \xnz.mem_r [816] = \xnz.mem_r_816_sv2v_reg ;
  assign \xnz.mem_r [815] = \xnz.mem_r_815_sv2v_reg ;
  assign \xnz.mem_r [814] = \xnz.mem_r_814_sv2v_reg ;
  assign \xnz.mem_r [813] = \xnz.mem_r_813_sv2v_reg ;
  assign \xnz.mem_r [812] = \xnz.mem_r_812_sv2v_reg ;
  assign \xnz.mem_r [811] = \xnz.mem_r_811_sv2v_reg ;
  assign \xnz.mem_r [810] = \xnz.mem_r_810_sv2v_reg ;
  assign \xnz.mem_r [809] = \xnz.mem_r_809_sv2v_reg ;
  assign \xnz.mem_r [808] = \xnz.mem_r_808_sv2v_reg ;
  assign \xnz.mem_r [807] = \xnz.mem_r_807_sv2v_reg ;
  assign \xnz.mem_r [806] = \xnz.mem_r_806_sv2v_reg ;
  assign \xnz.mem_r [805] = \xnz.mem_r_805_sv2v_reg ;
  assign \xnz.mem_r [804] = \xnz.mem_r_804_sv2v_reg ;
  assign \xnz.mem_r [803] = \xnz.mem_r_803_sv2v_reg ;
  assign \xnz.mem_r [802] = \xnz.mem_r_802_sv2v_reg ;
  assign \xnz.mem_r [801] = \xnz.mem_r_801_sv2v_reg ;
  assign \xnz.mem_r [800] = \xnz.mem_r_800_sv2v_reg ;
  assign \xnz.mem_r [799] = \xnz.mem_r_799_sv2v_reg ;
  assign \xnz.mem_r [798] = \xnz.mem_r_798_sv2v_reg ;
  assign \xnz.mem_r [797] = \xnz.mem_r_797_sv2v_reg ;
  assign \xnz.mem_r [796] = \xnz.mem_r_796_sv2v_reg ;
  assign \xnz.mem_r [795] = \xnz.mem_r_795_sv2v_reg ;
  assign \xnz.mem_r [794] = \xnz.mem_r_794_sv2v_reg ;
  assign \xnz.mem_r [793] = \xnz.mem_r_793_sv2v_reg ;
  assign \xnz.mem_r [792] = \xnz.mem_r_792_sv2v_reg ;
  assign \xnz.mem_r [791] = \xnz.mem_r_791_sv2v_reg ;
  assign \xnz.mem_r [790] = \xnz.mem_r_790_sv2v_reg ;
  assign \xnz.mem_r [789] = \xnz.mem_r_789_sv2v_reg ;
  assign \xnz.mem_r [788] = \xnz.mem_r_788_sv2v_reg ;
  assign \xnz.mem_r [787] = \xnz.mem_r_787_sv2v_reg ;
  assign \xnz.mem_r [786] = \xnz.mem_r_786_sv2v_reg ;
  assign \xnz.mem_r [785] = \xnz.mem_r_785_sv2v_reg ;
  assign \xnz.mem_r [784] = \xnz.mem_r_784_sv2v_reg ;
  assign \xnz.mem_r [783] = \xnz.mem_r_783_sv2v_reg ;
  assign \xnz.mem_r [782] = \xnz.mem_r_782_sv2v_reg ;
  assign \xnz.mem_r [781] = \xnz.mem_r_781_sv2v_reg ;
  assign \xnz.mem_r [780] = \xnz.mem_r_780_sv2v_reg ;
  assign \xnz.mem_r [779] = \xnz.mem_r_779_sv2v_reg ;
  assign \xnz.mem_r [778] = \xnz.mem_r_778_sv2v_reg ;
  assign \xnz.mem_r [777] = \xnz.mem_r_777_sv2v_reg ;
  assign \xnz.mem_r [776] = \xnz.mem_r_776_sv2v_reg ;
  assign \xnz.mem_r [775] = \xnz.mem_r_775_sv2v_reg ;
  assign \xnz.mem_r [774] = \xnz.mem_r_774_sv2v_reg ;
  assign \xnz.mem_r [773] = \xnz.mem_r_773_sv2v_reg ;
  assign \xnz.mem_r [772] = \xnz.mem_r_772_sv2v_reg ;
  assign \xnz.mem_r [771] = \xnz.mem_r_771_sv2v_reg ;
  assign \xnz.mem_r [770] = \xnz.mem_r_770_sv2v_reg ;
  assign \xnz.mem_r [769] = \xnz.mem_r_769_sv2v_reg ;
  assign \xnz.mem_r [768] = \xnz.mem_r_768_sv2v_reg ;
  assign \xnz.mem_r [767] = \xnz.mem_r_767_sv2v_reg ;
  assign \xnz.mem_r [766] = \xnz.mem_r_766_sv2v_reg ;
  assign \xnz.mem_r [765] = \xnz.mem_r_765_sv2v_reg ;
  assign \xnz.mem_r [764] = \xnz.mem_r_764_sv2v_reg ;
  assign \xnz.mem_r [763] = \xnz.mem_r_763_sv2v_reg ;
  assign \xnz.mem_r [762] = \xnz.mem_r_762_sv2v_reg ;
  assign \xnz.mem_r [761] = \xnz.mem_r_761_sv2v_reg ;
  assign \xnz.mem_r [760] = \xnz.mem_r_760_sv2v_reg ;
  assign \xnz.mem_r [759] = \xnz.mem_r_759_sv2v_reg ;
  assign \xnz.mem_r [758] = \xnz.mem_r_758_sv2v_reg ;
  assign \xnz.mem_r [757] = \xnz.mem_r_757_sv2v_reg ;
  assign \xnz.mem_r [756] = \xnz.mem_r_756_sv2v_reg ;
  assign \xnz.mem_r [755] = \xnz.mem_r_755_sv2v_reg ;
  assign \xnz.mem_r [754] = \xnz.mem_r_754_sv2v_reg ;
  assign \xnz.mem_r [753] = \xnz.mem_r_753_sv2v_reg ;
  assign \xnz.mem_r [752] = \xnz.mem_r_752_sv2v_reg ;
  assign \xnz.mem_r [751] = \xnz.mem_r_751_sv2v_reg ;
  assign \xnz.mem_r [750] = \xnz.mem_r_750_sv2v_reg ;
  assign \xnz.mem_r [749] = \xnz.mem_r_749_sv2v_reg ;
  assign \xnz.mem_r [748] = \xnz.mem_r_748_sv2v_reg ;
  assign \xnz.mem_r [747] = \xnz.mem_r_747_sv2v_reg ;
  assign \xnz.mem_r [746] = \xnz.mem_r_746_sv2v_reg ;
  assign \xnz.mem_r [745] = \xnz.mem_r_745_sv2v_reg ;
  assign \xnz.mem_r [744] = \xnz.mem_r_744_sv2v_reg ;
  assign \xnz.mem_r [743] = \xnz.mem_r_743_sv2v_reg ;
  assign \xnz.mem_r [742] = \xnz.mem_r_742_sv2v_reg ;
  assign \xnz.mem_r [741] = \xnz.mem_r_741_sv2v_reg ;
  assign \xnz.mem_r [740] = \xnz.mem_r_740_sv2v_reg ;
  assign \xnz.mem_r [739] = \xnz.mem_r_739_sv2v_reg ;
  assign \xnz.mem_r [738] = \xnz.mem_r_738_sv2v_reg ;
  assign \xnz.mem_r [737] = \xnz.mem_r_737_sv2v_reg ;
  assign \xnz.mem_r [736] = \xnz.mem_r_736_sv2v_reg ;
  assign \xnz.mem_r [735] = \xnz.mem_r_735_sv2v_reg ;
  assign \xnz.mem_r [734] = \xnz.mem_r_734_sv2v_reg ;
  assign \xnz.mem_r [733] = \xnz.mem_r_733_sv2v_reg ;
  assign \xnz.mem_r [732] = \xnz.mem_r_732_sv2v_reg ;
  assign \xnz.mem_r [731] = \xnz.mem_r_731_sv2v_reg ;
  assign \xnz.mem_r [730] = \xnz.mem_r_730_sv2v_reg ;
  assign \xnz.mem_r [729] = \xnz.mem_r_729_sv2v_reg ;
  assign \xnz.mem_r [728] = \xnz.mem_r_728_sv2v_reg ;
  assign \xnz.mem_r [727] = \xnz.mem_r_727_sv2v_reg ;
  assign \xnz.mem_r [726] = \xnz.mem_r_726_sv2v_reg ;
  assign \xnz.mem_r [725] = \xnz.mem_r_725_sv2v_reg ;
  assign \xnz.mem_r [724] = \xnz.mem_r_724_sv2v_reg ;
  assign \xnz.mem_r [723] = \xnz.mem_r_723_sv2v_reg ;
  assign \xnz.mem_r [722] = \xnz.mem_r_722_sv2v_reg ;
  assign \xnz.mem_r [721] = \xnz.mem_r_721_sv2v_reg ;
  assign \xnz.mem_r [720] = \xnz.mem_r_720_sv2v_reg ;
  assign \xnz.mem_r [719] = \xnz.mem_r_719_sv2v_reg ;
  assign \xnz.mem_r [718] = \xnz.mem_r_718_sv2v_reg ;
  assign \xnz.mem_r [717] = \xnz.mem_r_717_sv2v_reg ;
  assign \xnz.mem_r [716] = \xnz.mem_r_716_sv2v_reg ;
  assign \xnz.mem_r [715] = \xnz.mem_r_715_sv2v_reg ;
  assign \xnz.mem_r [714] = \xnz.mem_r_714_sv2v_reg ;
  assign \xnz.mem_r [713] = \xnz.mem_r_713_sv2v_reg ;
  assign \xnz.mem_r [712] = \xnz.mem_r_712_sv2v_reg ;
  assign \xnz.mem_r [711] = \xnz.mem_r_711_sv2v_reg ;
  assign \xnz.mem_r [710] = \xnz.mem_r_710_sv2v_reg ;
  assign \xnz.mem_r [709] = \xnz.mem_r_709_sv2v_reg ;
  assign \xnz.mem_r [708] = \xnz.mem_r_708_sv2v_reg ;
  assign \xnz.mem_r [707] = \xnz.mem_r_707_sv2v_reg ;
  assign \xnz.mem_r [706] = \xnz.mem_r_706_sv2v_reg ;
  assign \xnz.mem_r [705] = \xnz.mem_r_705_sv2v_reg ;
  assign \xnz.mem_r [704] = \xnz.mem_r_704_sv2v_reg ;
  assign \xnz.mem_r [703] = \xnz.mem_r_703_sv2v_reg ;
  assign \xnz.mem_r [702] = \xnz.mem_r_702_sv2v_reg ;
  assign \xnz.mem_r [701] = \xnz.mem_r_701_sv2v_reg ;
  assign \xnz.mem_r [700] = \xnz.mem_r_700_sv2v_reg ;
  assign \xnz.mem_r [699] = \xnz.mem_r_699_sv2v_reg ;
  assign \xnz.mem_r [698] = \xnz.mem_r_698_sv2v_reg ;
  assign \xnz.mem_r [697] = \xnz.mem_r_697_sv2v_reg ;
  assign \xnz.mem_r [696] = \xnz.mem_r_696_sv2v_reg ;
  assign \xnz.mem_r [695] = \xnz.mem_r_695_sv2v_reg ;
  assign \xnz.mem_r [694] = \xnz.mem_r_694_sv2v_reg ;
  assign \xnz.mem_r [693] = \xnz.mem_r_693_sv2v_reg ;
  assign \xnz.mem_r [692] = \xnz.mem_r_692_sv2v_reg ;
  assign \xnz.mem_r [691] = \xnz.mem_r_691_sv2v_reg ;
  assign \xnz.mem_r [690] = \xnz.mem_r_690_sv2v_reg ;
  assign \xnz.mem_r [689] = \xnz.mem_r_689_sv2v_reg ;
  assign \xnz.mem_r [688] = \xnz.mem_r_688_sv2v_reg ;
  assign \xnz.mem_r [687] = \xnz.mem_r_687_sv2v_reg ;
  assign \xnz.mem_r [686] = \xnz.mem_r_686_sv2v_reg ;
  assign \xnz.mem_r [685] = \xnz.mem_r_685_sv2v_reg ;
  assign \xnz.mem_r [684] = \xnz.mem_r_684_sv2v_reg ;
  assign \xnz.mem_r [683] = \xnz.mem_r_683_sv2v_reg ;
  assign \xnz.mem_r [682] = \xnz.mem_r_682_sv2v_reg ;
  assign \xnz.mem_r [681] = \xnz.mem_r_681_sv2v_reg ;
  assign \xnz.mem_r [680] = \xnz.mem_r_680_sv2v_reg ;
  assign \xnz.mem_r [679] = \xnz.mem_r_679_sv2v_reg ;
  assign \xnz.mem_r [678] = \xnz.mem_r_678_sv2v_reg ;
  assign \xnz.mem_r [677] = \xnz.mem_r_677_sv2v_reg ;
  assign \xnz.mem_r [676] = \xnz.mem_r_676_sv2v_reg ;
  assign \xnz.mem_r [675] = \xnz.mem_r_675_sv2v_reg ;
  assign \xnz.mem_r [674] = \xnz.mem_r_674_sv2v_reg ;
  assign \xnz.mem_r [673] = \xnz.mem_r_673_sv2v_reg ;
  assign \xnz.mem_r [672] = \xnz.mem_r_672_sv2v_reg ;
  assign \xnz.mem_r [671] = \xnz.mem_r_671_sv2v_reg ;
  assign \xnz.mem_r [670] = \xnz.mem_r_670_sv2v_reg ;
  assign \xnz.mem_r [669] = \xnz.mem_r_669_sv2v_reg ;
  assign \xnz.mem_r [668] = \xnz.mem_r_668_sv2v_reg ;
  assign \xnz.mem_r [667] = \xnz.mem_r_667_sv2v_reg ;
  assign \xnz.mem_r [666] = \xnz.mem_r_666_sv2v_reg ;
  assign \xnz.mem_r [665] = \xnz.mem_r_665_sv2v_reg ;
  assign \xnz.mem_r [664] = \xnz.mem_r_664_sv2v_reg ;
  assign \xnz.mem_r [663] = \xnz.mem_r_663_sv2v_reg ;
  assign \xnz.mem_r [662] = \xnz.mem_r_662_sv2v_reg ;
  assign \xnz.mem_r [661] = \xnz.mem_r_661_sv2v_reg ;
  assign \xnz.mem_r [660] = \xnz.mem_r_660_sv2v_reg ;
  assign \xnz.mem_r [659] = \xnz.mem_r_659_sv2v_reg ;
  assign \xnz.mem_r [658] = \xnz.mem_r_658_sv2v_reg ;
  assign \xnz.mem_r [657] = \xnz.mem_r_657_sv2v_reg ;
  assign \xnz.mem_r [656] = \xnz.mem_r_656_sv2v_reg ;
  assign \xnz.mem_r [655] = \xnz.mem_r_655_sv2v_reg ;
  assign \xnz.mem_r [654] = \xnz.mem_r_654_sv2v_reg ;
  assign \xnz.mem_r [653] = \xnz.mem_r_653_sv2v_reg ;
  assign \xnz.mem_r [652] = \xnz.mem_r_652_sv2v_reg ;
  assign \xnz.mem_r [651] = \xnz.mem_r_651_sv2v_reg ;
  assign \xnz.mem_r [650] = \xnz.mem_r_650_sv2v_reg ;
  assign \xnz.mem_r [649] = \xnz.mem_r_649_sv2v_reg ;
  assign \xnz.mem_r [648] = \xnz.mem_r_648_sv2v_reg ;
  assign \xnz.mem_r [647] = \xnz.mem_r_647_sv2v_reg ;
  assign \xnz.mem_r [646] = \xnz.mem_r_646_sv2v_reg ;
  assign \xnz.mem_r [645] = \xnz.mem_r_645_sv2v_reg ;
  assign \xnz.mem_r [644] = \xnz.mem_r_644_sv2v_reg ;
  assign \xnz.mem_r [643] = \xnz.mem_r_643_sv2v_reg ;
  assign \xnz.mem_r [642] = \xnz.mem_r_642_sv2v_reg ;
  assign \xnz.mem_r [641] = \xnz.mem_r_641_sv2v_reg ;
  assign \xnz.mem_r [640] = \xnz.mem_r_640_sv2v_reg ;
  assign \xnz.mem_r [639] = \xnz.mem_r_639_sv2v_reg ;
  assign \xnz.mem_r [638] = \xnz.mem_r_638_sv2v_reg ;
  assign \xnz.mem_r [637] = \xnz.mem_r_637_sv2v_reg ;
  assign \xnz.mem_r [636] = \xnz.mem_r_636_sv2v_reg ;
  assign \xnz.mem_r [635] = \xnz.mem_r_635_sv2v_reg ;
  assign \xnz.mem_r [634] = \xnz.mem_r_634_sv2v_reg ;
  assign \xnz.mem_r [633] = \xnz.mem_r_633_sv2v_reg ;
  assign \xnz.mem_r [632] = \xnz.mem_r_632_sv2v_reg ;
  assign \xnz.mem_r [631] = \xnz.mem_r_631_sv2v_reg ;
  assign \xnz.mem_r [630] = \xnz.mem_r_630_sv2v_reg ;
  assign \xnz.mem_r [629] = \xnz.mem_r_629_sv2v_reg ;
  assign \xnz.mem_r [628] = \xnz.mem_r_628_sv2v_reg ;
  assign \xnz.mem_r [627] = \xnz.mem_r_627_sv2v_reg ;
  assign \xnz.mem_r [626] = \xnz.mem_r_626_sv2v_reg ;
  assign \xnz.mem_r [625] = \xnz.mem_r_625_sv2v_reg ;
  assign \xnz.mem_r [624] = \xnz.mem_r_624_sv2v_reg ;
  assign \xnz.mem_r [623] = \xnz.mem_r_623_sv2v_reg ;
  assign \xnz.mem_r [622] = \xnz.mem_r_622_sv2v_reg ;
  assign \xnz.mem_r [621] = \xnz.mem_r_621_sv2v_reg ;
  assign \xnz.mem_r [620] = \xnz.mem_r_620_sv2v_reg ;
  assign \xnz.mem_r [619] = \xnz.mem_r_619_sv2v_reg ;
  assign \xnz.mem_r [618] = \xnz.mem_r_618_sv2v_reg ;
  assign \xnz.mem_r [617] = \xnz.mem_r_617_sv2v_reg ;
  assign \xnz.mem_r [616] = \xnz.mem_r_616_sv2v_reg ;
  assign \xnz.mem_r [615] = \xnz.mem_r_615_sv2v_reg ;
  assign \xnz.mem_r [614] = \xnz.mem_r_614_sv2v_reg ;
  assign \xnz.mem_r [613] = \xnz.mem_r_613_sv2v_reg ;
  assign \xnz.mem_r [612] = \xnz.mem_r_612_sv2v_reg ;
  assign \xnz.mem_r [611] = \xnz.mem_r_611_sv2v_reg ;
  assign \xnz.mem_r [610] = \xnz.mem_r_610_sv2v_reg ;
  assign \xnz.mem_r [609] = \xnz.mem_r_609_sv2v_reg ;
  assign \xnz.mem_r [608] = \xnz.mem_r_608_sv2v_reg ;
  assign \xnz.mem_r [607] = \xnz.mem_r_607_sv2v_reg ;
  assign \xnz.mem_r [606] = \xnz.mem_r_606_sv2v_reg ;
  assign \xnz.mem_r [605] = \xnz.mem_r_605_sv2v_reg ;
  assign \xnz.mem_r [604] = \xnz.mem_r_604_sv2v_reg ;
  assign \xnz.mem_r [603] = \xnz.mem_r_603_sv2v_reg ;
  assign \xnz.mem_r [602] = \xnz.mem_r_602_sv2v_reg ;
  assign \xnz.mem_r [601] = \xnz.mem_r_601_sv2v_reg ;
  assign \xnz.mem_r [600] = \xnz.mem_r_600_sv2v_reg ;
  assign \xnz.mem_r [599] = \xnz.mem_r_599_sv2v_reg ;
  assign \xnz.mem_r [598] = \xnz.mem_r_598_sv2v_reg ;
  assign \xnz.mem_r [597] = \xnz.mem_r_597_sv2v_reg ;
  assign \xnz.mem_r [596] = \xnz.mem_r_596_sv2v_reg ;
  assign \xnz.mem_r [595] = \xnz.mem_r_595_sv2v_reg ;
  assign \xnz.mem_r [594] = \xnz.mem_r_594_sv2v_reg ;
  assign \xnz.mem_r [593] = \xnz.mem_r_593_sv2v_reg ;
  assign \xnz.mem_r [592] = \xnz.mem_r_592_sv2v_reg ;
  assign \xnz.mem_r [591] = \xnz.mem_r_591_sv2v_reg ;
  assign \xnz.mem_r [590] = \xnz.mem_r_590_sv2v_reg ;
  assign \xnz.mem_r [589] = \xnz.mem_r_589_sv2v_reg ;
  assign \xnz.mem_r [588] = \xnz.mem_r_588_sv2v_reg ;
  assign \xnz.mem_r [587] = \xnz.mem_r_587_sv2v_reg ;
  assign \xnz.mem_r [586] = \xnz.mem_r_586_sv2v_reg ;
  assign \xnz.mem_r [585] = \xnz.mem_r_585_sv2v_reg ;
  assign \xnz.mem_r [584] = \xnz.mem_r_584_sv2v_reg ;
  assign \xnz.mem_r [583] = \xnz.mem_r_583_sv2v_reg ;
  assign \xnz.mem_r [582] = \xnz.mem_r_582_sv2v_reg ;
  assign \xnz.mem_r [581] = \xnz.mem_r_581_sv2v_reg ;
  assign \xnz.mem_r [580] = \xnz.mem_r_580_sv2v_reg ;
  assign \xnz.mem_r [579] = \xnz.mem_r_579_sv2v_reg ;
  assign \xnz.mem_r [578] = \xnz.mem_r_578_sv2v_reg ;
  assign \xnz.mem_r [577] = \xnz.mem_r_577_sv2v_reg ;
  assign \xnz.mem_r [576] = \xnz.mem_r_576_sv2v_reg ;
  assign \xnz.mem_r [575] = \xnz.mem_r_575_sv2v_reg ;
  assign \xnz.mem_r [574] = \xnz.mem_r_574_sv2v_reg ;
  assign \xnz.mem_r [573] = \xnz.mem_r_573_sv2v_reg ;
  assign \xnz.mem_r [572] = \xnz.mem_r_572_sv2v_reg ;
  assign \xnz.mem_r [571] = \xnz.mem_r_571_sv2v_reg ;
  assign \xnz.mem_r [570] = \xnz.mem_r_570_sv2v_reg ;
  assign \xnz.mem_r [569] = \xnz.mem_r_569_sv2v_reg ;
  assign \xnz.mem_r [568] = \xnz.mem_r_568_sv2v_reg ;
  assign \xnz.mem_r [567] = \xnz.mem_r_567_sv2v_reg ;
  assign \xnz.mem_r [566] = \xnz.mem_r_566_sv2v_reg ;
  assign \xnz.mem_r [565] = \xnz.mem_r_565_sv2v_reg ;
  assign \xnz.mem_r [564] = \xnz.mem_r_564_sv2v_reg ;
  assign \xnz.mem_r [563] = \xnz.mem_r_563_sv2v_reg ;
  assign \xnz.mem_r [562] = \xnz.mem_r_562_sv2v_reg ;
  assign \xnz.mem_r [561] = \xnz.mem_r_561_sv2v_reg ;
  assign \xnz.mem_r [560] = \xnz.mem_r_560_sv2v_reg ;
  assign \xnz.mem_r [559] = \xnz.mem_r_559_sv2v_reg ;
  assign \xnz.mem_r [558] = \xnz.mem_r_558_sv2v_reg ;
  assign \xnz.mem_r [557] = \xnz.mem_r_557_sv2v_reg ;
  assign \xnz.mem_r [556] = \xnz.mem_r_556_sv2v_reg ;
  assign \xnz.mem_r [555] = \xnz.mem_r_555_sv2v_reg ;
  assign \xnz.mem_r [554] = \xnz.mem_r_554_sv2v_reg ;
  assign \xnz.mem_r [553] = \xnz.mem_r_553_sv2v_reg ;
  assign \xnz.mem_r [552] = \xnz.mem_r_552_sv2v_reg ;
  assign \xnz.mem_r [551] = \xnz.mem_r_551_sv2v_reg ;
  assign \xnz.mem_r [550] = \xnz.mem_r_550_sv2v_reg ;
  assign \xnz.mem_r [549] = \xnz.mem_r_549_sv2v_reg ;
  assign \xnz.mem_r [548] = \xnz.mem_r_548_sv2v_reg ;
  assign \xnz.mem_r [547] = \xnz.mem_r_547_sv2v_reg ;
  assign \xnz.mem_r [546] = \xnz.mem_r_546_sv2v_reg ;
  assign \xnz.mem_r [545] = \xnz.mem_r_545_sv2v_reg ;
  assign \xnz.mem_r [544] = \xnz.mem_r_544_sv2v_reg ;
  assign \xnz.mem_r [543] = \xnz.mem_r_543_sv2v_reg ;
  assign \xnz.mem_r [542] = \xnz.mem_r_542_sv2v_reg ;
  assign \xnz.mem_r [541] = \xnz.mem_r_541_sv2v_reg ;
  assign \xnz.mem_r [540] = \xnz.mem_r_540_sv2v_reg ;
  assign \xnz.mem_r [539] = \xnz.mem_r_539_sv2v_reg ;
  assign \xnz.mem_r [538] = \xnz.mem_r_538_sv2v_reg ;
  assign \xnz.mem_r [537] = \xnz.mem_r_537_sv2v_reg ;
  assign \xnz.mem_r [536] = \xnz.mem_r_536_sv2v_reg ;
  assign \xnz.mem_r [535] = \xnz.mem_r_535_sv2v_reg ;
  assign \xnz.mem_r [534] = \xnz.mem_r_534_sv2v_reg ;
  assign \xnz.mem_r [533] = \xnz.mem_r_533_sv2v_reg ;
  assign \xnz.mem_r [532] = \xnz.mem_r_532_sv2v_reg ;
  assign \xnz.mem_r [531] = \xnz.mem_r_531_sv2v_reg ;
  assign \xnz.mem_r [530] = \xnz.mem_r_530_sv2v_reg ;
  assign \xnz.mem_r [529] = \xnz.mem_r_529_sv2v_reg ;
  assign \xnz.mem_r [528] = \xnz.mem_r_528_sv2v_reg ;
  assign \xnz.mem_r [527] = \xnz.mem_r_527_sv2v_reg ;
  assign \xnz.mem_r [526] = \xnz.mem_r_526_sv2v_reg ;
  assign \xnz.mem_r [525] = \xnz.mem_r_525_sv2v_reg ;
  assign \xnz.mem_r [524] = \xnz.mem_r_524_sv2v_reg ;
  assign \xnz.mem_r [523] = \xnz.mem_r_523_sv2v_reg ;
  assign \xnz.mem_r [522] = \xnz.mem_r_522_sv2v_reg ;
  assign \xnz.mem_r [521] = \xnz.mem_r_521_sv2v_reg ;
  assign \xnz.mem_r [520] = \xnz.mem_r_520_sv2v_reg ;
  assign \xnz.mem_r [519] = \xnz.mem_r_519_sv2v_reg ;
  assign \xnz.mem_r [518] = \xnz.mem_r_518_sv2v_reg ;
  assign \xnz.mem_r [517] = \xnz.mem_r_517_sv2v_reg ;
  assign \xnz.mem_r [516] = \xnz.mem_r_516_sv2v_reg ;
  assign \xnz.mem_r [515] = \xnz.mem_r_515_sv2v_reg ;
  assign \xnz.mem_r [514] = \xnz.mem_r_514_sv2v_reg ;
  assign \xnz.mem_r [513] = \xnz.mem_r_513_sv2v_reg ;
  assign \xnz.mem_r [512] = \xnz.mem_r_512_sv2v_reg ;
  assign \xnz.mem_r [511] = \xnz.mem_r_511_sv2v_reg ;
  assign \xnz.mem_r [510] = \xnz.mem_r_510_sv2v_reg ;
  assign \xnz.mem_r [509] = \xnz.mem_r_509_sv2v_reg ;
  assign \xnz.mem_r [508] = \xnz.mem_r_508_sv2v_reg ;
  assign \xnz.mem_r [507] = \xnz.mem_r_507_sv2v_reg ;
  assign \xnz.mem_r [506] = \xnz.mem_r_506_sv2v_reg ;
  assign \xnz.mem_r [505] = \xnz.mem_r_505_sv2v_reg ;
  assign \xnz.mem_r [504] = \xnz.mem_r_504_sv2v_reg ;
  assign \xnz.mem_r [503] = \xnz.mem_r_503_sv2v_reg ;
  assign \xnz.mem_r [502] = \xnz.mem_r_502_sv2v_reg ;
  assign \xnz.mem_r [501] = \xnz.mem_r_501_sv2v_reg ;
  assign \xnz.mem_r [500] = \xnz.mem_r_500_sv2v_reg ;
  assign \xnz.mem_r [499] = \xnz.mem_r_499_sv2v_reg ;
  assign \xnz.mem_r [498] = \xnz.mem_r_498_sv2v_reg ;
  assign \xnz.mem_r [497] = \xnz.mem_r_497_sv2v_reg ;
  assign \xnz.mem_r [496] = \xnz.mem_r_496_sv2v_reg ;
  assign \xnz.mem_r [495] = \xnz.mem_r_495_sv2v_reg ;
  assign \xnz.mem_r [494] = \xnz.mem_r_494_sv2v_reg ;
  assign \xnz.mem_r [493] = \xnz.mem_r_493_sv2v_reg ;
  assign \xnz.mem_r [492] = \xnz.mem_r_492_sv2v_reg ;
  assign \xnz.mem_r [491] = \xnz.mem_r_491_sv2v_reg ;
  assign \xnz.mem_r [490] = \xnz.mem_r_490_sv2v_reg ;
  assign \xnz.mem_r [489] = \xnz.mem_r_489_sv2v_reg ;
  assign \xnz.mem_r [488] = \xnz.mem_r_488_sv2v_reg ;
  assign \xnz.mem_r [487] = \xnz.mem_r_487_sv2v_reg ;
  assign \xnz.mem_r [486] = \xnz.mem_r_486_sv2v_reg ;
  assign \xnz.mem_r [485] = \xnz.mem_r_485_sv2v_reg ;
  assign \xnz.mem_r [484] = \xnz.mem_r_484_sv2v_reg ;
  assign \xnz.mem_r [483] = \xnz.mem_r_483_sv2v_reg ;
  assign \xnz.mem_r [482] = \xnz.mem_r_482_sv2v_reg ;
  assign \xnz.mem_r [481] = \xnz.mem_r_481_sv2v_reg ;
  assign \xnz.mem_r [480] = \xnz.mem_r_480_sv2v_reg ;
  assign \xnz.mem_r [479] = \xnz.mem_r_479_sv2v_reg ;
  assign \xnz.mem_r [478] = \xnz.mem_r_478_sv2v_reg ;
  assign \xnz.mem_r [477] = \xnz.mem_r_477_sv2v_reg ;
  assign \xnz.mem_r [476] = \xnz.mem_r_476_sv2v_reg ;
  assign \xnz.mem_r [475] = \xnz.mem_r_475_sv2v_reg ;
  assign \xnz.mem_r [474] = \xnz.mem_r_474_sv2v_reg ;
  assign \xnz.mem_r [473] = \xnz.mem_r_473_sv2v_reg ;
  assign \xnz.mem_r [472] = \xnz.mem_r_472_sv2v_reg ;
  assign \xnz.mem_r [471] = \xnz.mem_r_471_sv2v_reg ;
  assign \xnz.mem_r [470] = \xnz.mem_r_470_sv2v_reg ;
  assign \xnz.mem_r [469] = \xnz.mem_r_469_sv2v_reg ;
  assign \xnz.mem_r [468] = \xnz.mem_r_468_sv2v_reg ;
  assign \xnz.mem_r [467] = \xnz.mem_r_467_sv2v_reg ;
  assign \xnz.mem_r [466] = \xnz.mem_r_466_sv2v_reg ;
  assign \xnz.mem_r [465] = \xnz.mem_r_465_sv2v_reg ;
  assign \xnz.mem_r [464] = \xnz.mem_r_464_sv2v_reg ;
  assign \xnz.mem_r [463] = \xnz.mem_r_463_sv2v_reg ;
  assign \xnz.mem_r [462] = \xnz.mem_r_462_sv2v_reg ;
  assign \xnz.mem_r [461] = \xnz.mem_r_461_sv2v_reg ;
  assign \xnz.mem_r [460] = \xnz.mem_r_460_sv2v_reg ;
  assign \xnz.mem_r [459] = \xnz.mem_r_459_sv2v_reg ;
  assign \xnz.mem_r [458] = \xnz.mem_r_458_sv2v_reg ;
  assign \xnz.mem_r [457] = \xnz.mem_r_457_sv2v_reg ;
  assign \xnz.mem_r [456] = \xnz.mem_r_456_sv2v_reg ;
  assign \xnz.mem_r [455] = \xnz.mem_r_455_sv2v_reg ;
  assign \xnz.mem_r [454] = \xnz.mem_r_454_sv2v_reg ;
  assign \xnz.mem_r [453] = \xnz.mem_r_453_sv2v_reg ;
  assign \xnz.mem_r [452] = \xnz.mem_r_452_sv2v_reg ;
  assign \xnz.mem_r [451] = \xnz.mem_r_451_sv2v_reg ;
  assign \xnz.mem_r [450] = \xnz.mem_r_450_sv2v_reg ;
  assign \xnz.mem_r [449] = \xnz.mem_r_449_sv2v_reg ;
  assign \xnz.mem_r [448] = \xnz.mem_r_448_sv2v_reg ;
  assign \xnz.mem_r [447] = \xnz.mem_r_447_sv2v_reg ;
  assign \xnz.mem_r [446] = \xnz.mem_r_446_sv2v_reg ;
  assign \xnz.mem_r [445] = \xnz.mem_r_445_sv2v_reg ;
  assign \xnz.mem_r [444] = \xnz.mem_r_444_sv2v_reg ;
  assign \xnz.mem_r [443] = \xnz.mem_r_443_sv2v_reg ;
  assign \xnz.mem_r [442] = \xnz.mem_r_442_sv2v_reg ;
  assign \xnz.mem_r [441] = \xnz.mem_r_441_sv2v_reg ;
  assign \xnz.mem_r [440] = \xnz.mem_r_440_sv2v_reg ;
  assign \xnz.mem_r [439] = \xnz.mem_r_439_sv2v_reg ;
  assign \xnz.mem_r [438] = \xnz.mem_r_438_sv2v_reg ;
  assign \xnz.mem_r [437] = \xnz.mem_r_437_sv2v_reg ;
  assign \xnz.mem_r [436] = \xnz.mem_r_436_sv2v_reg ;
  assign \xnz.mem_r [435] = \xnz.mem_r_435_sv2v_reg ;
  assign \xnz.mem_r [434] = \xnz.mem_r_434_sv2v_reg ;
  assign \xnz.mem_r [433] = \xnz.mem_r_433_sv2v_reg ;
  assign \xnz.mem_r [432] = \xnz.mem_r_432_sv2v_reg ;
  assign \xnz.mem_r [431] = \xnz.mem_r_431_sv2v_reg ;
  assign \xnz.mem_r [430] = \xnz.mem_r_430_sv2v_reg ;
  assign \xnz.mem_r [429] = \xnz.mem_r_429_sv2v_reg ;
  assign \xnz.mem_r [428] = \xnz.mem_r_428_sv2v_reg ;
  assign \xnz.mem_r [427] = \xnz.mem_r_427_sv2v_reg ;
  assign \xnz.mem_r [426] = \xnz.mem_r_426_sv2v_reg ;
  assign \xnz.mem_r [425] = \xnz.mem_r_425_sv2v_reg ;
  assign \xnz.mem_r [424] = \xnz.mem_r_424_sv2v_reg ;
  assign \xnz.mem_r [423] = \xnz.mem_r_423_sv2v_reg ;
  assign \xnz.mem_r [422] = \xnz.mem_r_422_sv2v_reg ;
  assign \xnz.mem_r [421] = \xnz.mem_r_421_sv2v_reg ;
  assign \xnz.mem_r [420] = \xnz.mem_r_420_sv2v_reg ;
  assign \xnz.mem_r [419] = \xnz.mem_r_419_sv2v_reg ;
  assign \xnz.mem_r [418] = \xnz.mem_r_418_sv2v_reg ;
  assign \xnz.mem_r [417] = \xnz.mem_r_417_sv2v_reg ;
  assign \xnz.mem_r [416] = \xnz.mem_r_416_sv2v_reg ;
  assign \xnz.mem_r [415] = \xnz.mem_r_415_sv2v_reg ;
  assign \xnz.mem_r [414] = \xnz.mem_r_414_sv2v_reg ;
  assign \xnz.mem_r [413] = \xnz.mem_r_413_sv2v_reg ;
  assign \xnz.mem_r [412] = \xnz.mem_r_412_sv2v_reg ;
  assign \xnz.mem_r [411] = \xnz.mem_r_411_sv2v_reg ;
  assign \xnz.mem_r [410] = \xnz.mem_r_410_sv2v_reg ;
  assign \xnz.mem_r [409] = \xnz.mem_r_409_sv2v_reg ;
  assign \xnz.mem_r [408] = \xnz.mem_r_408_sv2v_reg ;
  assign \xnz.mem_r [407] = \xnz.mem_r_407_sv2v_reg ;
  assign \xnz.mem_r [406] = \xnz.mem_r_406_sv2v_reg ;
  assign \xnz.mem_r [405] = \xnz.mem_r_405_sv2v_reg ;
  assign \xnz.mem_r [404] = \xnz.mem_r_404_sv2v_reg ;
  assign \xnz.mem_r [403] = \xnz.mem_r_403_sv2v_reg ;
  assign \xnz.mem_r [402] = \xnz.mem_r_402_sv2v_reg ;
  assign \xnz.mem_r [401] = \xnz.mem_r_401_sv2v_reg ;
  assign \xnz.mem_r [400] = \xnz.mem_r_400_sv2v_reg ;
  assign \xnz.mem_r [399] = \xnz.mem_r_399_sv2v_reg ;
  assign \xnz.mem_r [398] = \xnz.mem_r_398_sv2v_reg ;
  assign \xnz.mem_r [397] = \xnz.mem_r_397_sv2v_reg ;
  assign \xnz.mem_r [396] = \xnz.mem_r_396_sv2v_reg ;
  assign \xnz.mem_r [395] = \xnz.mem_r_395_sv2v_reg ;
  assign \xnz.mem_r [394] = \xnz.mem_r_394_sv2v_reg ;
  assign \xnz.mem_r [393] = \xnz.mem_r_393_sv2v_reg ;
  assign \xnz.mem_r [392] = \xnz.mem_r_392_sv2v_reg ;
  assign \xnz.mem_r [391] = \xnz.mem_r_391_sv2v_reg ;
  assign \xnz.mem_r [390] = \xnz.mem_r_390_sv2v_reg ;
  assign \xnz.mem_r [389] = \xnz.mem_r_389_sv2v_reg ;
  assign \xnz.mem_r [388] = \xnz.mem_r_388_sv2v_reg ;
  assign \xnz.mem_r [387] = \xnz.mem_r_387_sv2v_reg ;
  assign \xnz.mem_r [386] = \xnz.mem_r_386_sv2v_reg ;
  assign \xnz.mem_r [385] = \xnz.mem_r_385_sv2v_reg ;
  assign \xnz.mem_r [384] = \xnz.mem_r_384_sv2v_reg ;
  assign \xnz.mem_r [383] = \xnz.mem_r_383_sv2v_reg ;
  assign \xnz.mem_r [382] = \xnz.mem_r_382_sv2v_reg ;
  assign \xnz.mem_r [381] = \xnz.mem_r_381_sv2v_reg ;
  assign \xnz.mem_r [380] = \xnz.mem_r_380_sv2v_reg ;
  assign \xnz.mem_r [379] = \xnz.mem_r_379_sv2v_reg ;
  assign \xnz.mem_r [378] = \xnz.mem_r_378_sv2v_reg ;
  assign \xnz.mem_r [377] = \xnz.mem_r_377_sv2v_reg ;
  assign \xnz.mem_r [376] = \xnz.mem_r_376_sv2v_reg ;
  assign \xnz.mem_r [375] = \xnz.mem_r_375_sv2v_reg ;
  assign \xnz.mem_r [374] = \xnz.mem_r_374_sv2v_reg ;
  assign \xnz.mem_r [373] = \xnz.mem_r_373_sv2v_reg ;
  assign \xnz.mem_r [372] = \xnz.mem_r_372_sv2v_reg ;
  assign \xnz.mem_r [371] = \xnz.mem_r_371_sv2v_reg ;
  assign \xnz.mem_r [370] = \xnz.mem_r_370_sv2v_reg ;
  assign \xnz.mem_r [369] = \xnz.mem_r_369_sv2v_reg ;
  assign \xnz.mem_r [368] = \xnz.mem_r_368_sv2v_reg ;
  assign \xnz.mem_r [367] = \xnz.mem_r_367_sv2v_reg ;
  assign \xnz.mem_r [366] = \xnz.mem_r_366_sv2v_reg ;
  assign \xnz.mem_r [365] = \xnz.mem_r_365_sv2v_reg ;
  assign \xnz.mem_r [364] = \xnz.mem_r_364_sv2v_reg ;
  assign \xnz.mem_r [363] = \xnz.mem_r_363_sv2v_reg ;
  assign \xnz.mem_r [362] = \xnz.mem_r_362_sv2v_reg ;
  assign \xnz.mem_r [361] = \xnz.mem_r_361_sv2v_reg ;
  assign \xnz.mem_r [360] = \xnz.mem_r_360_sv2v_reg ;
  assign \xnz.mem_r [359] = \xnz.mem_r_359_sv2v_reg ;
  assign \xnz.mem_r [358] = \xnz.mem_r_358_sv2v_reg ;
  assign \xnz.mem_r [357] = \xnz.mem_r_357_sv2v_reg ;
  assign \xnz.mem_r [356] = \xnz.mem_r_356_sv2v_reg ;
  assign \xnz.mem_r [355] = \xnz.mem_r_355_sv2v_reg ;
  assign \xnz.mem_r [354] = \xnz.mem_r_354_sv2v_reg ;
  assign \xnz.mem_r [353] = \xnz.mem_r_353_sv2v_reg ;
  assign \xnz.mem_r [352] = \xnz.mem_r_352_sv2v_reg ;
  assign \xnz.mem_r [351] = \xnz.mem_r_351_sv2v_reg ;
  assign \xnz.mem_r [350] = \xnz.mem_r_350_sv2v_reg ;
  assign \xnz.mem_r [349] = \xnz.mem_r_349_sv2v_reg ;
  assign \xnz.mem_r [348] = \xnz.mem_r_348_sv2v_reg ;
  assign \xnz.mem_r [347] = \xnz.mem_r_347_sv2v_reg ;
  assign \xnz.mem_r [346] = \xnz.mem_r_346_sv2v_reg ;
  assign \xnz.mem_r [345] = \xnz.mem_r_345_sv2v_reg ;
  assign \xnz.mem_r [344] = \xnz.mem_r_344_sv2v_reg ;
  assign \xnz.mem_r [343] = \xnz.mem_r_343_sv2v_reg ;
  assign \xnz.mem_r [342] = \xnz.mem_r_342_sv2v_reg ;
  assign \xnz.mem_r [341] = \xnz.mem_r_341_sv2v_reg ;
  assign \xnz.mem_r [340] = \xnz.mem_r_340_sv2v_reg ;
  assign \xnz.mem_r [339] = \xnz.mem_r_339_sv2v_reg ;
  assign \xnz.mem_r [338] = \xnz.mem_r_338_sv2v_reg ;
  assign \xnz.mem_r [337] = \xnz.mem_r_337_sv2v_reg ;
  assign \xnz.mem_r [336] = \xnz.mem_r_336_sv2v_reg ;
  assign \xnz.mem_r [335] = \xnz.mem_r_335_sv2v_reg ;
  assign \xnz.mem_r [334] = \xnz.mem_r_334_sv2v_reg ;
  assign \xnz.mem_r [333] = \xnz.mem_r_333_sv2v_reg ;
  assign \xnz.mem_r [332] = \xnz.mem_r_332_sv2v_reg ;
  assign \xnz.mem_r [331] = \xnz.mem_r_331_sv2v_reg ;
  assign \xnz.mem_r [330] = \xnz.mem_r_330_sv2v_reg ;
  assign \xnz.mem_r [329] = \xnz.mem_r_329_sv2v_reg ;
  assign \xnz.mem_r [328] = \xnz.mem_r_328_sv2v_reg ;
  assign \xnz.mem_r [327] = \xnz.mem_r_327_sv2v_reg ;
  assign \xnz.mem_r [326] = \xnz.mem_r_326_sv2v_reg ;
  assign \xnz.mem_r [325] = \xnz.mem_r_325_sv2v_reg ;
  assign \xnz.mem_r [324] = \xnz.mem_r_324_sv2v_reg ;
  assign \xnz.mem_r [323] = \xnz.mem_r_323_sv2v_reg ;
  assign \xnz.mem_r [322] = \xnz.mem_r_322_sv2v_reg ;
  assign \xnz.mem_r [321] = \xnz.mem_r_321_sv2v_reg ;
  assign \xnz.mem_r [320] = \xnz.mem_r_320_sv2v_reg ;
  assign \xnz.mem_r [319] = \xnz.mem_r_319_sv2v_reg ;
  assign \xnz.mem_r [318] = \xnz.mem_r_318_sv2v_reg ;
  assign \xnz.mem_r [317] = \xnz.mem_r_317_sv2v_reg ;
  assign \xnz.mem_r [316] = \xnz.mem_r_316_sv2v_reg ;
  assign \xnz.mem_r [315] = \xnz.mem_r_315_sv2v_reg ;
  assign \xnz.mem_r [314] = \xnz.mem_r_314_sv2v_reg ;
  assign \xnz.mem_r [313] = \xnz.mem_r_313_sv2v_reg ;
  assign \xnz.mem_r [312] = \xnz.mem_r_312_sv2v_reg ;
  assign \xnz.mem_r [311] = \xnz.mem_r_311_sv2v_reg ;
  assign \xnz.mem_r [310] = \xnz.mem_r_310_sv2v_reg ;
  assign \xnz.mem_r [309] = \xnz.mem_r_309_sv2v_reg ;
  assign \xnz.mem_r [308] = \xnz.mem_r_308_sv2v_reg ;
  assign \xnz.mem_r [307] = \xnz.mem_r_307_sv2v_reg ;
  assign \xnz.mem_r [306] = \xnz.mem_r_306_sv2v_reg ;
  assign \xnz.mem_r [305] = \xnz.mem_r_305_sv2v_reg ;
  assign \xnz.mem_r [304] = \xnz.mem_r_304_sv2v_reg ;
  assign \xnz.mem_r [303] = \xnz.mem_r_303_sv2v_reg ;
  assign \xnz.mem_r [302] = \xnz.mem_r_302_sv2v_reg ;
  assign \xnz.mem_r [301] = \xnz.mem_r_301_sv2v_reg ;
  assign \xnz.mem_r [300] = \xnz.mem_r_300_sv2v_reg ;
  assign \xnz.mem_r [299] = \xnz.mem_r_299_sv2v_reg ;
  assign \xnz.mem_r [298] = \xnz.mem_r_298_sv2v_reg ;
  assign \xnz.mem_r [297] = \xnz.mem_r_297_sv2v_reg ;
  assign \xnz.mem_r [296] = \xnz.mem_r_296_sv2v_reg ;
  assign \xnz.mem_r [295] = \xnz.mem_r_295_sv2v_reg ;
  assign \xnz.mem_r [294] = \xnz.mem_r_294_sv2v_reg ;
  assign \xnz.mem_r [293] = \xnz.mem_r_293_sv2v_reg ;
  assign \xnz.mem_r [292] = \xnz.mem_r_292_sv2v_reg ;
  assign \xnz.mem_r [291] = \xnz.mem_r_291_sv2v_reg ;
  assign \xnz.mem_r [290] = \xnz.mem_r_290_sv2v_reg ;
  assign \xnz.mem_r [289] = \xnz.mem_r_289_sv2v_reg ;
  assign \xnz.mem_r [288] = \xnz.mem_r_288_sv2v_reg ;
  assign \xnz.mem_r [287] = \xnz.mem_r_287_sv2v_reg ;
  assign \xnz.mem_r [286] = \xnz.mem_r_286_sv2v_reg ;
  assign \xnz.mem_r [285] = \xnz.mem_r_285_sv2v_reg ;
  assign \xnz.mem_r [284] = \xnz.mem_r_284_sv2v_reg ;
  assign \xnz.mem_r [283] = \xnz.mem_r_283_sv2v_reg ;
  assign \xnz.mem_r [282] = \xnz.mem_r_282_sv2v_reg ;
  assign \xnz.mem_r [281] = \xnz.mem_r_281_sv2v_reg ;
  assign \xnz.mem_r [280] = \xnz.mem_r_280_sv2v_reg ;
  assign \xnz.mem_r [279] = \xnz.mem_r_279_sv2v_reg ;
  assign \xnz.mem_r [278] = \xnz.mem_r_278_sv2v_reg ;
  assign \xnz.mem_r [277] = \xnz.mem_r_277_sv2v_reg ;
  assign \xnz.mem_r [276] = \xnz.mem_r_276_sv2v_reg ;
  assign \xnz.mem_r [275] = \xnz.mem_r_275_sv2v_reg ;
  assign \xnz.mem_r [274] = \xnz.mem_r_274_sv2v_reg ;
  assign \xnz.mem_r [273] = \xnz.mem_r_273_sv2v_reg ;
  assign \xnz.mem_r [272] = \xnz.mem_r_272_sv2v_reg ;
  assign \xnz.mem_r [271] = \xnz.mem_r_271_sv2v_reg ;
  assign \xnz.mem_r [270] = \xnz.mem_r_270_sv2v_reg ;
  assign \xnz.mem_r [269] = \xnz.mem_r_269_sv2v_reg ;
  assign \xnz.mem_r [268] = \xnz.mem_r_268_sv2v_reg ;
  assign \xnz.mem_r [267] = \xnz.mem_r_267_sv2v_reg ;
  assign \xnz.mem_r [266] = \xnz.mem_r_266_sv2v_reg ;
  assign \xnz.mem_r [265] = \xnz.mem_r_265_sv2v_reg ;
  assign \xnz.mem_r [264] = \xnz.mem_r_264_sv2v_reg ;
  assign \xnz.mem_r [263] = \xnz.mem_r_263_sv2v_reg ;
  assign \xnz.mem_r [262] = \xnz.mem_r_262_sv2v_reg ;
  assign \xnz.mem_r [261] = \xnz.mem_r_261_sv2v_reg ;
  assign \xnz.mem_r [260] = \xnz.mem_r_260_sv2v_reg ;
  assign \xnz.mem_r [259] = \xnz.mem_r_259_sv2v_reg ;
  assign \xnz.mem_r [258] = \xnz.mem_r_258_sv2v_reg ;
  assign \xnz.mem_r [257] = \xnz.mem_r_257_sv2v_reg ;
  assign \xnz.mem_r [256] = \xnz.mem_r_256_sv2v_reg ;
  assign \xnz.mem_r [255] = \xnz.mem_r_255_sv2v_reg ;
  assign \xnz.mem_r [254] = \xnz.mem_r_254_sv2v_reg ;
  assign \xnz.mem_r [253] = \xnz.mem_r_253_sv2v_reg ;
  assign \xnz.mem_r [252] = \xnz.mem_r_252_sv2v_reg ;
  assign \xnz.mem_r [251] = \xnz.mem_r_251_sv2v_reg ;
  assign \xnz.mem_r [250] = \xnz.mem_r_250_sv2v_reg ;
  assign \xnz.mem_r [249] = \xnz.mem_r_249_sv2v_reg ;
  assign \xnz.mem_r [248] = \xnz.mem_r_248_sv2v_reg ;
  assign \xnz.mem_r [247] = \xnz.mem_r_247_sv2v_reg ;
  assign \xnz.mem_r [246] = \xnz.mem_r_246_sv2v_reg ;
  assign \xnz.mem_r [245] = \xnz.mem_r_245_sv2v_reg ;
  assign \xnz.mem_r [244] = \xnz.mem_r_244_sv2v_reg ;
  assign \xnz.mem_r [243] = \xnz.mem_r_243_sv2v_reg ;
  assign \xnz.mem_r [242] = \xnz.mem_r_242_sv2v_reg ;
  assign \xnz.mem_r [241] = \xnz.mem_r_241_sv2v_reg ;
  assign \xnz.mem_r [240] = \xnz.mem_r_240_sv2v_reg ;
  assign \xnz.mem_r [239] = \xnz.mem_r_239_sv2v_reg ;
  assign \xnz.mem_r [238] = \xnz.mem_r_238_sv2v_reg ;
  assign \xnz.mem_r [237] = \xnz.mem_r_237_sv2v_reg ;
  assign \xnz.mem_r [236] = \xnz.mem_r_236_sv2v_reg ;
  assign \xnz.mem_r [235] = \xnz.mem_r_235_sv2v_reg ;
  assign \xnz.mem_r [234] = \xnz.mem_r_234_sv2v_reg ;
  assign \xnz.mem_r [233] = \xnz.mem_r_233_sv2v_reg ;
  assign \xnz.mem_r [232] = \xnz.mem_r_232_sv2v_reg ;
  assign \xnz.mem_r [231] = \xnz.mem_r_231_sv2v_reg ;
  assign \xnz.mem_r [230] = \xnz.mem_r_230_sv2v_reg ;
  assign \xnz.mem_r [229] = \xnz.mem_r_229_sv2v_reg ;
  assign \xnz.mem_r [228] = \xnz.mem_r_228_sv2v_reg ;
  assign \xnz.mem_r [227] = \xnz.mem_r_227_sv2v_reg ;
  assign \xnz.mem_r [226] = \xnz.mem_r_226_sv2v_reg ;
  assign \xnz.mem_r [225] = \xnz.mem_r_225_sv2v_reg ;
  assign \xnz.mem_r [224] = \xnz.mem_r_224_sv2v_reg ;
  assign \xnz.mem_r [223] = \xnz.mem_r_223_sv2v_reg ;
  assign \xnz.mem_r [222] = \xnz.mem_r_222_sv2v_reg ;
  assign \xnz.mem_r [221] = \xnz.mem_r_221_sv2v_reg ;
  assign \xnz.mem_r [220] = \xnz.mem_r_220_sv2v_reg ;
  assign \xnz.mem_r [219] = \xnz.mem_r_219_sv2v_reg ;
  assign \xnz.mem_r [218] = \xnz.mem_r_218_sv2v_reg ;
  assign \xnz.mem_r [217] = \xnz.mem_r_217_sv2v_reg ;
  assign \xnz.mem_r [216] = \xnz.mem_r_216_sv2v_reg ;
  assign \xnz.mem_r [215] = \xnz.mem_r_215_sv2v_reg ;
  assign \xnz.mem_r [214] = \xnz.mem_r_214_sv2v_reg ;
  assign \xnz.mem_r [213] = \xnz.mem_r_213_sv2v_reg ;
  assign \xnz.mem_r [212] = \xnz.mem_r_212_sv2v_reg ;
  assign \xnz.mem_r [211] = \xnz.mem_r_211_sv2v_reg ;
  assign \xnz.mem_r [210] = \xnz.mem_r_210_sv2v_reg ;
  assign \xnz.mem_r [209] = \xnz.mem_r_209_sv2v_reg ;
  assign \xnz.mem_r [208] = \xnz.mem_r_208_sv2v_reg ;
  assign \xnz.mem_r [207] = \xnz.mem_r_207_sv2v_reg ;
  assign \xnz.mem_r [206] = \xnz.mem_r_206_sv2v_reg ;
  assign \xnz.mem_r [205] = \xnz.mem_r_205_sv2v_reg ;
  assign \xnz.mem_r [204] = \xnz.mem_r_204_sv2v_reg ;
  assign \xnz.mem_r [203] = \xnz.mem_r_203_sv2v_reg ;
  assign \xnz.mem_r [202] = \xnz.mem_r_202_sv2v_reg ;
  assign \xnz.mem_r [201] = \xnz.mem_r_201_sv2v_reg ;
  assign \xnz.mem_r [200] = \xnz.mem_r_200_sv2v_reg ;
  assign \xnz.mem_r [199] = \xnz.mem_r_199_sv2v_reg ;
  assign \xnz.mem_r [198] = \xnz.mem_r_198_sv2v_reg ;
  assign \xnz.mem_r [197] = \xnz.mem_r_197_sv2v_reg ;
  assign \xnz.mem_r [196] = \xnz.mem_r_196_sv2v_reg ;
  assign \xnz.mem_r [195] = \xnz.mem_r_195_sv2v_reg ;
  assign \xnz.mem_r [194] = \xnz.mem_r_194_sv2v_reg ;
  assign \xnz.mem_r [193] = \xnz.mem_r_193_sv2v_reg ;
  assign \xnz.mem_r [192] = \xnz.mem_r_192_sv2v_reg ;
  assign \xnz.mem_r [191] = \xnz.mem_r_191_sv2v_reg ;
  assign \xnz.mem_r [190] = \xnz.mem_r_190_sv2v_reg ;
  assign \xnz.mem_r [189] = \xnz.mem_r_189_sv2v_reg ;
  assign \xnz.mem_r [188] = \xnz.mem_r_188_sv2v_reg ;
  assign \xnz.mem_r [187] = \xnz.mem_r_187_sv2v_reg ;
  assign \xnz.mem_r [186] = \xnz.mem_r_186_sv2v_reg ;
  assign \xnz.mem_r [185] = \xnz.mem_r_185_sv2v_reg ;
  assign \xnz.mem_r [184] = \xnz.mem_r_184_sv2v_reg ;
  assign \xnz.mem_r [183] = \xnz.mem_r_183_sv2v_reg ;
  assign \xnz.mem_r [182] = \xnz.mem_r_182_sv2v_reg ;
  assign \xnz.mem_r [181] = \xnz.mem_r_181_sv2v_reg ;
  assign \xnz.mem_r [180] = \xnz.mem_r_180_sv2v_reg ;
  assign \xnz.mem_r [179] = \xnz.mem_r_179_sv2v_reg ;
  assign \xnz.mem_r [178] = \xnz.mem_r_178_sv2v_reg ;
  assign \xnz.mem_r [177] = \xnz.mem_r_177_sv2v_reg ;
  assign \xnz.mem_r [176] = \xnz.mem_r_176_sv2v_reg ;
  assign \xnz.mem_r [175] = \xnz.mem_r_175_sv2v_reg ;
  assign \xnz.mem_r [174] = \xnz.mem_r_174_sv2v_reg ;
  assign \xnz.mem_r [173] = \xnz.mem_r_173_sv2v_reg ;
  assign \xnz.mem_r [172] = \xnz.mem_r_172_sv2v_reg ;
  assign \xnz.mem_r [171] = \xnz.mem_r_171_sv2v_reg ;
  assign \xnz.mem_r [170] = \xnz.mem_r_170_sv2v_reg ;
  assign \xnz.mem_r [169] = \xnz.mem_r_169_sv2v_reg ;
  assign \xnz.mem_r [168] = \xnz.mem_r_168_sv2v_reg ;
  assign \xnz.mem_r [167] = \xnz.mem_r_167_sv2v_reg ;
  assign \xnz.mem_r [166] = \xnz.mem_r_166_sv2v_reg ;
  assign \xnz.mem_r [165] = \xnz.mem_r_165_sv2v_reg ;
  assign \xnz.mem_r [164] = \xnz.mem_r_164_sv2v_reg ;
  assign \xnz.mem_r [163] = \xnz.mem_r_163_sv2v_reg ;
  assign \xnz.mem_r [162] = \xnz.mem_r_162_sv2v_reg ;
  assign \xnz.mem_r [161] = \xnz.mem_r_161_sv2v_reg ;
  assign \xnz.mem_r [160] = \xnz.mem_r_160_sv2v_reg ;
  assign \xnz.mem_r [159] = \xnz.mem_r_159_sv2v_reg ;
  assign \xnz.mem_r [158] = \xnz.mem_r_158_sv2v_reg ;
  assign \xnz.mem_r [157] = \xnz.mem_r_157_sv2v_reg ;
  assign \xnz.mem_r [156] = \xnz.mem_r_156_sv2v_reg ;
  assign \xnz.mem_r [155] = \xnz.mem_r_155_sv2v_reg ;
  assign \xnz.mem_r [154] = \xnz.mem_r_154_sv2v_reg ;
  assign \xnz.mem_r [153] = \xnz.mem_r_153_sv2v_reg ;
  assign \xnz.mem_r [152] = \xnz.mem_r_152_sv2v_reg ;
  assign \xnz.mem_r [151] = \xnz.mem_r_151_sv2v_reg ;
  assign \xnz.mem_r [150] = \xnz.mem_r_150_sv2v_reg ;
  assign \xnz.mem_r [149] = \xnz.mem_r_149_sv2v_reg ;
  assign \xnz.mem_r [148] = \xnz.mem_r_148_sv2v_reg ;
  assign \xnz.mem_r [147] = \xnz.mem_r_147_sv2v_reg ;
  assign \xnz.mem_r [146] = \xnz.mem_r_146_sv2v_reg ;
  assign \xnz.mem_r [145] = \xnz.mem_r_145_sv2v_reg ;
  assign \xnz.mem_r [144] = \xnz.mem_r_144_sv2v_reg ;
  assign \xnz.mem_r [143] = \xnz.mem_r_143_sv2v_reg ;
  assign \xnz.mem_r [142] = \xnz.mem_r_142_sv2v_reg ;
  assign \xnz.mem_r [141] = \xnz.mem_r_141_sv2v_reg ;
  assign \xnz.mem_r [140] = \xnz.mem_r_140_sv2v_reg ;
  assign \xnz.mem_r [139] = \xnz.mem_r_139_sv2v_reg ;
  assign \xnz.mem_r [138] = \xnz.mem_r_138_sv2v_reg ;
  assign \xnz.mem_r [137] = \xnz.mem_r_137_sv2v_reg ;
  assign \xnz.mem_r [136] = \xnz.mem_r_136_sv2v_reg ;
  assign \xnz.mem_r [135] = \xnz.mem_r_135_sv2v_reg ;
  assign \xnz.mem_r [134] = \xnz.mem_r_134_sv2v_reg ;
  assign \xnz.mem_r [133] = \xnz.mem_r_133_sv2v_reg ;
  assign \xnz.mem_r [132] = \xnz.mem_r_132_sv2v_reg ;
  assign \xnz.mem_r [131] = \xnz.mem_r_131_sv2v_reg ;
  assign \xnz.mem_r [130] = \xnz.mem_r_130_sv2v_reg ;
  assign \xnz.mem_r [129] = \xnz.mem_r_129_sv2v_reg ;
  assign \xnz.mem_r [128] = \xnz.mem_r_128_sv2v_reg ;
  assign \xnz.mem_r [127] = \xnz.mem_r_127_sv2v_reg ;
  assign \xnz.mem_r [126] = \xnz.mem_r_126_sv2v_reg ;
  assign \xnz.mem_r [125] = \xnz.mem_r_125_sv2v_reg ;
  assign \xnz.mem_r [124] = \xnz.mem_r_124_sv2v_reg ;
  assign \xnz.mem_r [123] = \xnz.mem_r_123_sv2v_reg ;
  assign \xnz.mem_r [122] = \xnz.mem_r_122_sv2v_reg ;
  assign \xnz.mem_r [121] = \xnz.mem_r_121_sv2v_reg ;
  assign \xnz.mem_r [120] = \xnz.mem_r_120_sv2v_reg ;
  assign \xnz.mem_r [119] = \xnz.mem_r_119_sv2v_reg ;
  assign \xnz.mem_r [118] = \xnz.mem_r_118_sv2v_reg ;
  assign \xnz.mem_r [117] = \xnz.mem_r_117_sv2v_reg ;
  assign \xnz.mem_r [116] = \xnz.mem_r_116_sv2v_reg ;
  assign \xnz.mem_r [115] = \xnz.mem_r_115_sv2v_reg ;
  assign \xnz.mem_r [114] = \xnz.mem_r_114_sv2v_reg ;
  assign \xnz.mem_r [113] = \xnz.mem_r_113_sv2v_reg ;
  assign \xnz.mem_r [112] = \xnz.mem_r_112_sv2v_reg ;
  assign \xnz.mem_r [111] = \xnz.mem_r_111_sv2v_reg ;
  assign \xnz.mem_r [110] = \xnz.mem_r_110_sv2v_reg ;
  assign \xnz.mem_r [109] = \xnz.mem_r_109_sv2v_reg ;
  assign \xnz.mem_r [108] = \xnz.mem_r_108_sv2v_reg ;
  assign \xnz.mem_r [107] = \xnz.mem_r_107_sv2v_reg ;
  assign \xnz.mem_r [106] = \xnz.mem_r_106_sv2v_reg ;
  assign \xnz.mem_r [105] = \xnz.mem_r_105_sv2v_reg ;
  assign \xnz.mem_r [104] = \xnz.mem_r_104_sv2v_reg ;
  assign \xnz.mem_r [103] = \xnz.mem_r_103_sv2v_reg ;
  assign \xnz.mem_r [102] = \xnz.mem_r_102_sv2v_reg ;
  assign \xnz.mem_r [101] = \xnz.mem_r_101_sv2v_reg ;
  assign \xnz.mem_r [100] = \xnz.mem_r_100_sv2v_reg ;
  assign \xnz.mem_r [99] = \xnz.mem_r_99_sv2v_reg ;
  assign \xnz.mem_r [98] = \xnz.mem_r_98_sv2v_reg ;
  assign \xnz.mem_r [97] = \xnz.mem_r_97_sv2v_reg ;
  assign \xnz.mem_r [96] = \xnz.mem_r_96_sv2v_reg ;
  assign \xnz.mem_r [95] = \xnz.mem_r_95_sv2v_reg ;
  assign \xnz.mem_r [94] = \xnz.mem_r_94_sv2v_reg ;
  assign \xnz.mem_r [93] = \xnz.mem_r_93_sv2v_reg ;
  assign \xnz.mem_r [92] = \xnz.mem_r_92_sv2v_reg ;
  assign \xnz.mem_r [91] = \xnz.mem_r_91_sv2v_reg ;
  assign \xnz.mem_r [90] = \xnz.mem_r_90_sv2v_reg ;
  assign \xnz.mem_r [89] = \xnz.mem_r_89_sv2v_reg ;
  assign \xnz.mem_r [88] = \xnz.mem_r_88_sv2v_reg ;
  assign \xnz.mem_r [87] = \xnz.mem_r_87_sv2v_reg ;
  assign \xnz.mem_r [86] = \xnz.mem_r_86_sv2v_reg ;
  assign \xnz.mem_r [85] = \xnz.mem_r_85_sv2v_reg ;
  assign \xnz.mem_r [84] = \xnz.mem_r_84_sv2v_reg ;
  assign \xnz.mem_r [83] = \xnz.mem_r_83_sv2v_reg ;
  assign \xnz.mem_r [82] = \xnz.mem_r_82_sv2v_reg ;
  assign \xnz.mem_r [81] = \xnz.mem_r_81_sv2v_reg ;
  assign \xnz.mem_r [80] = \xnz.mem_r_80_sv2v_reg ;
  assign \xnz.mem_r [79] = \xnz.mem_r_79_sv2v_reg ;
  assign \xnz.mem_r [78] = \xnz.mem_r_78_sv2v_reg ;
  assign \xnz.mem_r [77] = \xnz.mem_r_77_sv2v_reg ;
  assign \xnz.mem_r [76] = \xnz.mem_r_76_sv2v_reg ;
  assign \xnz.mem_r [75] = \xnz.mem_r_75_sv2v_reg ;
  assign \xnz.mem_r [74] = \xnz.mem_r_74_sv2v_reg ;
  assign \xnz.mem_r [73] = \xnz.mem_r_73_sv2v_reg ;
  assign \xnz.mem_r [72] = \xnz.mem_r_72_sv2v_reg ;
  assign \xnz.mem_r [71] = \xnz.mem_r_71_sv2v_reg ;
  assign \xnz.mem_r [70] = \xnz.mem_r_70_sv2v_reg ;
  assign \xnz.mem_r [69] = \xnz.mem_r_69_sv2v_reg ;
  assign \xnz.mem_r [68] = \xnz.mem_r_68_sv2v_reg ;
  assign \xnz.mem_r [67] = \xnz.mem_r_67_sv2v_reg ;
  assign \xnz.mem_r [66] = \xnz.mem_r_66_sv2v_reg ;
  assign \xnz.mem_r [65] = \xnz.mem_r_65_sv2v_reg ;
  assign \xnz.mem_r [64] = \xnz.mem_r_64_sv2v_reg ;
  assign \xnz.mem_r [63] = \xnz.mem_r_63_sv2v_reg ;
  assign \xnz.mem_r [62] = \xnz.mem_r_62_sv2v_reg ;
  assign \xnz.mem_r [61] = \xnz.mem_r_61_sv2v_reg ;
  assign \xnz.mem_r [60] = \xnz.mem_r_60_sv2v_reg ;
  assign \xnz.mem_r [59] = \xnz.mem_r_59_sv2v_reg ;
  assign \xnz.mem_r [58] = \xnz.mem_r_58_sv2v_reg ;
  assign \xnz.mem_r [57] = \xnz.mem_r_57_sv2v_reg ;
  assign \xnz.mem_r [56] = \xnz.mem_r_56_sv2v_reg ;
  assign \xnz.mem_r [55] = \xnz.mem_r_55_sv2v_reg ;
  assign \xnz.mem_r [54] = \xnz.mem_r_54_sv2v_reg ;
  assign \xnz.mem_r [53] = \xnz.mem_r_53_sv2v_reg ;
  assign \xnz.mem_r [52] = \xnz.mem_r_52_sv2v_reg ;
  assign \xnz.mem_r [51] = \xnz.mem_r_51_sv2v_reg ;
  assign \xnz.mem_r [50] = \xnz.mem_r_50_sv2v_reg ;
  assign \xnz.mem_r [49] = \xnz.mem_r_49_sv2v_reg ;
  assign \xnz.mem_r [48] = \xnz.mem_r_48_sv2v_reg ;
  assign \xnz.mem_r [47] = \xnz.mem_r_47_sv2v_reg ;
  assign \xnz.mem_r [46] = \xnz.mem_r_46_sv2v_reg ;
  assign \xnz.mem_r [45] = \xnz.mem_r_45_sv2v_reg ;
  assign \xnz.mem_r [44] = \xnz.mem_r_44_sv2v_reg ;
  assign \xnz.mem_r [43] = \xnz.mem_r_43_sv2v_reg ;
  assign \xnz.mem_r [42] = \xnz.mem_r_42_sv2v_reg ;
  assign \xnz.mem_r [41] = \xnz.mem_r_41_sv2v_reg ;
  assign \xnz.mem_r [40] = \xnz.mem_r_40_sv2v_reg ;
  assign \xnz.mem_r [39] = \xnz.mem_r_39_sv2v_reg ;
  assign \xnz.mem_r [38] = \xnz.mem_r_38_sv2v_reg ;
  assign \xnz.mem_r [37] = \xnz.mem_r_37_sv2v_reg ;
  assign \xnz.mem_r [36] = \xnz.mem_r_36_sv2v_reg ;
  assign \xnz.mem_r [35] = \xnz.mem_r_35_sv2v_reg ;
  assign \xnz.mem_r [34] = \xnz.mem_r_34_sv2v_reg ;
  assign \xnz.mem_r [33] = \xnz.mem_r_33_sv2v_reg ;
  assign \xnz.mem_r [32] = \xnz.mem_r_32_sv2v_reg ;
  assign \xnz.mem_r [31] = \xnz.mem_r_31_sv2v_reg ;
  assign \xnz.mem_r [30] = \xnz.mem_r_30_sv2v_reg ;
  assign \xnz.mem_r [29] = \xnz.mem_r_29_sv2v_reg ;
  assign \xnz.mem_r [28] = \xnz.mem_r_28_sv2v_reg ;
  assign \xnz.mem_r [27] = \xnz.mem_r_27_sv2v_reg ;
  assign \xnz.mem_r [26] = \xnz.mem_r_26_sv2v_reg ;
  assign \xnz.mem_r [25] = \xnz.mem_r_25_sv2v_reg ;
  assign \xnz.mem_r [24] = \xnz.mem_r_24_sv2v_reg ;
  assign \xnz.mem_r [23] = \xnz.mem_r_23_sv2v_reg ;
  assign \xnz.mem_r [22] = \xnz.mem_r_22_sv2v_reg ;
  assign \xnz.mem_r [21] = \xnz.mem_r_21_sv2v_reg ;
  assign \xnz.mem_r [20] = \xnz.mem_r_20_sv2v_reg ;
  assign \xnz.mem_r [19] = \xnz.mem_r_19_sv2v_reg ;
  assign \xnz.mem_r [18] = \xnz.mem_r_18_sv2v_reg ;
  assign \xnz.mem_r [17] = \xnz.mem_r_17_sv2v_reg ;
  assign \xnz.mem_r [16] = \xnz.mem_r_16_sv2v_reg ;
  assign \xnz.mem_r [15] = \xnz.mem_r_15_sv2v_reg ;
  assign \xnz.mem_r [14] = \xnz.mem_r_14_sv2v_reg ;
  assign \xnz.mem_r [13] = \xnz.mem_r_13_sv2v_reg ;
  assign \xnz.mem_r [12] = \xnz.mem_r_12_sv2v_reg ;
  assign \xnz.mem_r [11] = \xnz.mem_r_11_sv2v_reg ;
  assign \xnz.mem_r [10] = \xnz.mem_r_10_sv2v_reg ;
  assign \xnz.mem_r [9] = \xnz.mem_r_9_sv2v_reg ;
  assign \xnz.mem_r [8] = \xnz.mem_r_8_sv2v_reg ;
  assign \xnz.mem_r [7] = \xnz.mem_r_7_sv2v_reg ;
  assign \xnz.mem_r [6] = \xnz.mem_r_6_sv2v_reg ;
  assign \xnz.mem_r [5] = \xnz.mem_r_5_sv2v_reg ;
  assign \xnz.mem_r [4] = \xnz.mem_r_4_sv2v_reg ;
  assign \xnz.mem_r [3] = \xnz.mem_r_3_sv2v_reg ;
  assign \xnz.mem_r [2] = \xnz.mem_r_2_sv2v_reg ;
  assign \xnz.mem_r [1] = \xnz.mem_r_1_sv2v_reg ;
  assign \xnz.mem_r [0] = \xnz.mem_r_0_sv2v_reg ;
  assign r_data_o[32] = (N43)? \xnz.mem_r [32] : 
                        (N45)? \xnz.mem_r [65] : 
                        (N47)? \xnz.mem_r [98] : 
                        (N49)? \xnz.mem_r [131] : 
                        (N51)? \xnz.mem_r [164] : 
                        (N53)? \xnz.mem_r [197] : 
                        (N55)? \xnz.mem_r [230] : 
                        (N57)? \xnz.mem_r [263] : 
                        (N59)? \xnz.mem_r [296] : 
                        (N61)? \xnz.mem_r [329] : 
                        (N63)? \xnz.mem_r [362] : 
                        (N65)? \xnz.mem_r [395] : 
                        (N67)? \xnz.mem_r [428] : 
                        (N69)? \xnz.mem_r [461] : 
                        (N71)? \xnz.mem_r [494] : 
                        (N73)? \xnz.mem_r [527] : 
                        (N44)? \xnz.mem_r [560] : 
                        (N46)? \xnz.mem_r [593] : 
                        (N48)? \xnz.mem_r [626] : 
                        (N50)? \xnz.mem_r [659] : 
                        (N52)? \xnz.mem_r [692] : 
                        (N54)? \xnz.mem_r [725] : 
                        (N56)? \xnz.mem_r [758] : 
                        (N58)? \xnz.mem_r [791] : 
                        (N60)? \xnz.mem_r [824] : 
                        (N62)? \xnz.mem_r [857] : 
                        (N64)? \xnz.mem_r [890] : 
                        (N66)? \xnz.mem_r [923] : 
                        (N68)? \xnz.mem_r [956] : 
                        (N70)? \xnz.mem_r [989] : 
                        (N72)? \xnz.mem_r [1022] : 
                        (N74)? \xnz.mem_r [1055] : 1'b0;
  assign r_data_o[31] = (N43)? \xnz.mem_r [31] : 
                        (N45)? \xnz.mem_r [64] : 
                        (N47)? \xnz.mem_r [97] : 
                        (N49)? \xnz.mem_r [130] : 
                        (N51)? \xnz.mem_r [163] : 
                        (N53)? \xnz.mem_r [196] : 
                        (N55)? \xnz.mem_r [229] : 
                        (N57)? \xnz.mem_r [262] : 
                        (N59)? \xnz.mem_r [295] : 
                        (N61)? \xnz.mem_r [328] : 
                        (N63)? \xnz.mem_r [361] : 
                        (N65)? \xnz.mem_r [394] : 
                        (N67)? \xnz.mem_r [427] : 
                        (N69)? \xnz.mem_r [460] : 
                        (N71)? \xnz.mem_r [493] : 
                        (N73)? \xnz.mem_r [526] : 
                        (N44)? \xnz.mem_r [559] : 
                        (N46)? \xnz.mem_r [592] : 
                        (N48)? \xnz.mem_r [625] : 
                        (N50)? \xnz.mem_r [658] : 
                        (N52)? \xnz.mem_r [691] : 
                        (N54)? \xnz.mem_r [724] : 
                        (N56)? \xnz.mem_r [757] : 
                        (N58)? \xnz.mem_r [790] : 
                        (N60)? \xnz.mem_r [823] : 
                        (N62)? \xnz.mem_r [856] : 
                        (N64)? \xnz.mem_r [889] : 
                        (N66)? \xnz.mem_r [922] : 
                        (N68)? \xnz.mem_r [955] : 
                        (N70)? \xnz.mem_r [988] : 
                        (N72)? \xnz.mem_r [1021] : 
                        (N74)? \xnz.mem_r [1054] : 1'b0;
  assign r_data_o[30] = (N43)? \xnz.mem_r [30] : 
                        (N45)? \xnz.mem_r [63] : 
                        (N47)? \xnz.mem_r [96] : 
                        (N49)? \xnz.mem_r [129] : 
                        (N51)? \xnz.mem_r [162] : 
                        (N53)? \xnz.mem_r [195] : 
                        (N55)? \xnz.mem_r [228] : 
                        (N57)? \xnz.mem_r [261] : 
                        (N59)? \xnz.mem_r [294] : 
                        (N61)? \xnz.mem_r [327] : 
                        (N63)? \xnz.mem_r [360] : 
                        (N65)? \xnz.mem_r [393] : 
                        (N67)? \xnz.mem_r [426] : 
                        (N69)? \xnz.mem_r [459] : 
                        (N71)? \xnz.mem_r [492] : 
                        (N73)? \xnz.mem_r [525] : 
                        (N44)? \xnz.mem_r [558] : 
                        (N46)? \xnz.mem_r [591] : 
                        (N48)? \xnz.mem_r [624] : 
                        (N50)? \xnz.mem_r [657] : 
                        (N52)? \xnz.mem_r [690] : 
                        (N54)? \xnz.mem_r [723] : 
                        (N56)? \xnz.mem_r [756] : 
                        (N58)? \xnz.mem_r [789] : 
                        (N60)? \xnz.mem_r [822] : 
                        (N62)? \xnz.mem_r [855] : 
                        (N64)? \xnz.mem_r [888] : 
                        (N66)? \xnz.mem_r [921] : 
                        (N68)? \xnz.mem_r [954] : 
                        (N70)? \xnz.mem_r [987] : 
                        (N72)? \xnz.mem_r [1020] : 
                        (N74)? \xnz.mem_r [1053] : 1'b0;
  assign r_data_o[29] = (N43)? \xnz.mem_r [29] : 
                        (N45)? \xnz.mem_r [62] : 
                        (N47)? \xnz.mem_r [95] : 
                        (N49)? \xnz.mem_r [128] : 
                        (N51)? \xnz.mem_r [161] : 
                        (N53)? \xnz.mem_r [194] : 
                        (N55)? \xnz.mem_r [227] : 
                        (N57)? \xnz.mem_r [260] : 
                        (N59)? \xnz.mem_r [293] : 
                        (N61)? \xnz.mem_r [326] : 
                        (N63)? \xnz.mem_r [359] : 
                        (N65)? \xnz.mem_r [392] : 
                        (N67)? \xnz.mem_r [425] : 
                        (N69)? \xnz.mem_r [458] : 
                        (N71)? \xnz.mem_r [491] : 
                        (N73)? \xnz.mem_r [524] : 
                        (N44)? \xnz.mem_r [557] : 
                        (N46)? \xnz.mem_r [590] : 
                        (N48)? \xnz.mem_r [623] : 
                        (N50)? \xnz.mem_r [656] : 
                        (N52)? \xnz.mem_r [689] : 
                        (N54)? \xnz.mem_r [722] : 
                        (N56)? \xnz.mem_r [755] : 
                        (N58)? \xnz.mem_r [788] : 
                        (N60)? \xnz.mem_r [821] : 
                        (N62)? \xnz.mem_r [854] : 
                        (N64)? \xnz.mem_r [887] : 
                        (N66)? \xnz.mem_r [920] : 
                        (N68)? \xnz.mem_r [953] : 
                        (N70)? \xnz.mem_r [986] : 
                        (N72)? \xnz.mem_r [1019] : 
                        (N74)? \xnz.mem_r [1052] : 1'b0;
  assign r_data_o[28] = (N43)? \xnz.mem_r [28] : 
                        (N45)? \xnz.mem_r [61] : 
                        (N47)? \xnz.mem_r [94] : 
                        (N49)? \xnz.mem_r [127] : 
                        (N51)? \xnz.mem_r [160] : 
                        (N53)? \xnz.mem_r [193] : 
                        (N55)? \xnz.mem_r [226] : 
                        (N57)? \xnz.mem_r [259] : 
                        (N59)? \xnz.mem_r [292] : 
                        (N61)? \xnz.mem_r [325] : 
                        (N63)? \xnz.mem_r [358] : 
                        (N65)? \xnz.mem_r [391] : 
                        (N67)? \xnz.mem_r [424] : 
                        (N69)? \xnz.mem_r [457] : 
                        (N71)? \xnz.mem_r [490] : 
                        (N73)? \xnz.mem_r [523] : 
                        (N44)? \xnz.mem_r [556] : 
                        (N46)? \xnz.mem_r [589] : 
                        (N48)? \xnz.mem_r [622] : 
                        (N50)? \xnz.mem_r [655] : 
                        (N52)? \xnz.mem_r [688] : 
                        (N54)? \xnz.mem_r [721] : 
                        (N56)? \xnz.mem_r [754] : 
                        (N58)? \xnz.mem_r [787] : 
                        (N60)? \xnz.mem_r [820] : 
                        (N62)? \xnz.mem_r [853] : 
                        (N64)? \xnz.mem_r [886] : 
                        (N66)? \xnz.mem_r [919] : 
                        (N68)? \xnz.mem_r [952] : 
                        (N70)? \xnz.mem_r [985] : 
                        (N72)? \xnz.mem_r [1018] : 
                        (N74)? \xnz.mem_r [1051] : 1'b0;
  assign r_data_o[27] = (N43)? \xnz.mem_r [27] : 
                        (N45)? \xnz.mem_r [60] : 
                        (N47)? \xnz.mem_r [93] : 
                        (N49)? \xnz.mem_r [126] : 
                        (N51)? \xnz.mem_r [159] : 
                        (N53)? \xnz.mem_r [192] : 
                        (N55)? \xnz.mem_r [225] : 
                        (N57)? \xnz.mem_r [258] : 
                        (N59)? \xnz.mem_r [291] : 
                        (N61)? \xnz.mem_r [324] : 
                        (N63)? \xnz.mem_r [357] : 
                        (N65)? \xnz.mem_r [390] : 
                        (N67)? \xnz.mem_r [423] : 
                        (N69)? \xnz.mem_r [456] : 
                        (N71)? \xnz.mem_r [489] : 
                        (N73)? \xnz.mem_r [522] : 
                        (N44)? \xnz.mem_r [555] : 
                        (N46)? \xnz.mem_r [588] : 
                        (N48)? \xnz.mem_r [621] : 
                        (N50)? \xnz.mem_r [654] : 
                        (N52)? \xnz.mem_r [687] : 
                        (N54)? \xnz.mem_r [720] : 
                        (N56)? \xnz.mem_r [753] : 
                        (N58)? \xnz.mem_r [786] : 
                        (N60)? \xnz.mem_r [819] : 
                        (N62)? \xnz.mem_r [852] : 
                        (N64)? \xnz.mem_r [885] : 
                        (N66)? \xnz.mem_r [918] : 
                        (N68)? \xnz.mem_r [951] : 
                        (N70)? \xnz.mem_r [984] : 
                        (N72)? \xnz.mem_r [1017] : 
                        (N74)? \xnz.mem_r [1050] : 1'b0;
  assign r_data_o[26] = (N43)? \xnz.mem_r [26] : 
                        (N45)? \xnz.mem_r [59] : 
                        (N47)? \xnz.mem_r [92] : 
                        (N49)? \xnz.mem_r [125] : 
                        (N51)? \xnz.mem_r [158] : 
                        (N53)? \xnz.mem_r [191] : 
                        (N55)? \xnz.mem_r [224] : 
                        (N57)? \xnz.mem_r [257] : 
                        (N59)? \xnz.mem_r [290] : 
                        (N61)? \xnz.mem_r [323] : 
                        (N63)? \xnz.mem_r [356] : 
                        (N65)? \xnz.mem_r [389] : 
                        (N67)? \xnz.mem_r [422] : 
                        (N69)? \xnz.mem_r [455] : 
                        (N71)? \xnz.mem_r [488] : 
                        (N73)? \xnz.mem_r [521] : 
                        (N44)? \xnz.mem_r [554] : 
                        (N46)? \xnz.mem_r [587] : 
                        (N48)? \xnz.mem_r [620] : 
                        (N50)? \xnz.mem_r [653] : 
                        (N52)? \xnz.mem_r [686] : 
                        (N54)? \xnz.mem_r [719] : 
                        (N56)? \xnz.mem_r [752] : 
                        (N58)? \xnz.mem_r [785] : 
                        (N60)? \xnz.mem_r [818] : 
                        (N62)? \xnz.mem_r [851] : 
                        (N64)? \xnz.mem_r [884] : 
                        (N66)? \xnz.mem_r [917] : 
                        (N68)? \xnz.mem_r [950] : 
                        (N70)? \xnz.mem_r [983] : 
                        (N72)? \xnz.mem_r [1016] : 
                        (N74)? \xnz.mem_r [1049] : 1'b0;
  assign r_data_o[25] = (N43)? \xnz.mem_r [25] : 
                        (N45)? \xnz.mem_r [58] : 
                        (N47)? \xnz.mem_r [91] : 
                        (N49)? \xnz.mem_r [124] : 
                        (N51)? \xnz.mem_r [157] : 
                        (N53)? \xnz.mem_r [190] : 
                        (N55)? \xnz.mem_r [223] : 
                        (N57)? \xnz.mem_r [256] : 
                        (N59)? \xnz.mem_r [289] : 
                        (N61)? \xnz.mem_r [322] : 
                        (N63)? \xnz.mem_r [355] : 
                        (N65)? \xnz.mem_r [388] : 
                        (N67)? \xnz.mem_r [421] : 
                        (N69)? \xnz.mem_r [454] : 
                        (N71)? \xnz.mem_r [487] : 
                        (N73)? \xnz.mem_r [520] : 
                        (N44)? \xnz.mem_r [553] : 
                        (N46)? \xnz.mem_r [586] : 
                        (N48)? \xnz.mem_r [619] : 
                        (N50)? \xnz.mem_r [652] : 
                        (N52)? \xnz.mem_r [685] : 
                        (N54)? \xnz.mem_r [718] : 
                        (N56)? \xnz.mem_r [751] : 
                        (N58)? \xnz.mem_r [784] : 
                        (N60)? \xnz.mem_r [817] : 
                        (N62)? \xnz.mem_r [850] : 
                        (N64)? \xnz.mem_r [883] : 
                        (N66)? \xnz.mem_r [916] : 
                        (N68)? \xnz.mem_r [949] : 
                        (N70)? \xnz.mem_r [982] : 
                        (N72)? \xnz.mem_r [1015] : 
                        (N74)? \xnz.mem_r [1048] : 1'b0;
  assign r_data_o[24] = (N43)? \xnz.mem_r [24] : 
                        (N45)? \xnz.mem_r [57] : 
                        (N47)? \xnz.mem_r [90] : 
                        (N49)? \xnz.mem_r [123] : 
                        (N51)? \xnz.mem_r [156] : 
                        (N53)? \xnz.mem_r [189] : 
                        (N55)? \xnz.mem_r [222] : 
                        (N57)? \xnz.mem_r [255] : 
                        (N59)? \xnz.mem_r [288] : 
                        (N61)? \xnz.mem_r [321] : 
                        (N63)? \xnz.mem_r [354] : 
                        (N65)? \xnz.mem_r [387] : 
                        (N67)? \xnz.mem_r [420] : 
                        (N69)? \xnz.mem_r [453] : 
                        (N71)? \xnz.mem_r [486] : 
                        (N73)? \xnz.mem_r [519] : 
                        (N44)? \xnz.mem_r [552] : 
                        (N46)? \xnz.mem_r [585] : 
                        (N48)? \xnz.mem_r [618] : 
                        (N50)? \xnz.mem_r [651] : 
                        (N52)? \xnz.mem_r [684] : 
                        (N54)? \xnz.mem_r [717] : 
                        (N56)? \xnz.mem_r [750] : 
                        (N58)? \xnz.mem_r [783] : 
                        (N60)? \xnz.mem_r [816] : 
                        (N62)? \xnz.mem_r [849] : 
                        (N64)? \xnz.mem_r [882] : 
                        (N66)? \xnz.mem_r [915] : 
                        (N68)? \xnz.mem_r [948] : 
                        (N70)? \xnz.mem_r [981] : 
                        (N72)? \xnz.mem_r [1014] : 
                        (N74)? \xnz.mem_r [1047] : 1'b0;
  assign r_data_o[23] = (N43)? \xnz.mem_r [23] : 
                        (N45)? \xnz.mem_r [56] : 
                        (N47)? \xnz.mem_r [89] : 
                        (N49)? \xnz.mem_r [122] : 
                        (N51)? \xnz.mem_r [155] : 
                        (N53)? \xnz.mem_r [188] : 
                        (N55)? \xnz.mem_r [221] : 
                        (N57)? \xnz.mem_r [254] : 
                        (N59)? \xnz.mem_r [287] : 
                        (N61)? \xnz.mem_r [320] : 
                        (N63)? \xnz.mem_r [353] : 
                        (N65)? \xnz.mem_r [386] : 
                        (N67)? \xnz.mem_r [419] : 
                        (N69)? \xnz.mem_r [452] : 
                        (N71)? \xnz.mem_r [485] : 
                        (N73)? \xnz.mem_r [518] : 
                        (N44)? \xnz.mem_r [551] : 
                        (N46)? \xnz.mem_r [584] : 
                        (N48)? \xnz.mem_r [617] : 
                        (N50)? \xnz.mem_r [650] : 
                        (N52)? \xnz.mem_r [683] : 
                        (N54)? \xnz.mem_r [716] : 
                        (N56)? \xnz.mem_r [749] : 
                        (N58)? \xnz.mem_r [782] : 
                        (N60)? \xnz.mem_r [815] : 
                        (N62)? \xnz.mem_r [848] : 
                        (N64)? \xnz.mem_r [881] : 
                        (N66)? \xnz.mem_r [914] : 
                        (N68)? \xnz.mem_r [947] : 
                        (N70)? \xnz.mem_r [980] : 
                        (N72)? \xnz.mem_r [1013] : 
                        (N74)? \xnz.mem_r [1046] : 1'b0;
  assign r_data_o[22] = (N43)? \xnz.mem_r [22] : 
                        (N45)? \xnz.mem_r [55] : 
                        (N47)? \xnz.mem_r [88] : 
                        (N49)? \xnz.mem_r [121] : 
                        (N51)? \xnz.mem_r [154] : 
                        (N53)? \xnz.mem_r [187] : 
                        (N55)? \xnz.mem_r [220] : 
                        (N57)? \xnz.mem_r [253] : 
                        (N59)? \xnz.mem_r [286] : 
                        (N61)? \xnz.mem_r [319] : 
                        (N63)? \xnz.mem_r [352] : 
                        (N65)? \xnz.mem_r [385] : 
                        (N67)? \xnz.mem_r [418] : 
                        (N69)? \xnz.mem_r [451] : 
                        (N71)? \xnz.mem_r [484] : 
                        (N73)? \xnz.mem_r [517] : 
                        (N44)? \xnz.mem_r [550] : 
                        (N46)? \xnz.mem_r [583] : 
                        (N48)? \xnz.mem_r [616] : 
                        (N50)? \xnz.mem_r [649] : 
                        (N52)? \xnz.mem_r [682] : 
                        (N54)? \xnz.mem_r [715] : 
                        (N56)? \xnz.mem_r [748] : 
                        (N58)? \xnz.mem_r [781] : 
                        (N60)? \xnz.mem_r [814] : 
                        (N62)? \xnz.mem_r [847] : 
                        (N64)? \xnz.mem_r [880] : 
                        (N66)? \xnz.mem_r [913] : 
                        (N68)? \xnz.mem_r [946] : 
                        (N70)? \xnz.mem_r [979] : 
                        (N72)? \xnz.mem_r [1012] : 
                        (N74)? \xnz.mem_r [1045] : 1'b0;
  assign r_data_o[21] = (N43)? \xnz.mem_r [21] : 
                        (N45)? \xnz.mem_r [54] : 
                        (N47)? \xnz.mem_r [87] : 
                        (N49)? \xnz.mem_r [120] : 
                        (N51)? \xnz.mem_r [153] : 
                        (N53)? \xnz.mem_r [186] : 
                        (N55)? \xnz.mem_r [219] : 
                        (N57)? \xnz.mem_r [252] : 
                        (N59)? \xnz.mem_r [285] : 
                        (N61)? \xnz.mem_r [318] : 
                        (N63)? \xnz.mem_r [351] : 
                        (N65)? \xnz.mem_r [384] : 
                        (N67)? \xnz.mem_r [417] : 
                        (N69)? \xnz.mem_r [450] : 
                        (N71)? \xnz.mem_r [483] : 
                        (N73)? \xnz.mem_r [516] : 
                        (N44)? \xnz.mem_r [549] : 
                        (N46)? \xnz.mem_r [582] : 
                        (N48)? \xnz.mem_r [615] : 
                        (N50)? \xnz.mem_r [648] : 
                        (N52)? \xnz.mem_r [681] : 
                        (N54)? \xnz.mem_r [714] : 
                        (N56)? \xnz.mem_r [747] : 
                        (N58)? \xnz.mem_r [780] : 
                        (N60)? \xnz.mem_r [813] : 
                        (N62)? \xnz.mem_r [846] : 
                        (N64)? \xnz.mem_r [879] : 
                        (N66)? \xnz.mem_r [912] : 
                        (N68)? \xnz.mem_r [945] : 
                        (N70)? \xnz.mem_r [978] : 
                        (N72)? \xnz.mem_r [1011] : 
                        (N74)? \xnz.mem_r [1044] : 1'b0;
  assign r_data_o[20] = (N43)? \xnz.mem_r [20] : 
                        (N45)? \xnz.mem_r [53] : 
                        (N47)? \xnz.mem_r [86] : 
                        (N49)? \xnz.mem_r [119] : 
                        (N51)? \xnz.mem_r [152] : 
                        (N53)? \xnz.mem_r [185] : 
                        (N55)? \xnz.mem_r [218] : 
                        (N57)? \xnz.mem_r [251] : 
                        (N59)? \xnz.mem_r [284] : 
                        (N61)? \xnz.mem_r [317] : 
                        (N63)? \xnz.mem_r [350] : 
                        (N65)? \xnz.mem_r [383] : 
                        (N67)? \xnz.mem_r [416] : 
                        (N69)? \xnz.mem_r [449] : 
                        (N71)? \xnz.mem_r [482] : 
                        (N73)? \xnz.mem_r [515] : 
                        (N44)? \xnz.mem_r [548] : 
                        (N46)? \xnz.mem_r [581] : 
                        (N48)? \xnz.mem_r [614] : 
                        (N50)? \xnz.mem_r [647] : 
                        (N52)? \xnz.mem_r [680] : 
                        (N54)? \xnz.mem_r [713] : 
                        (N56)? \xnz.mem_r [746] : 
                        (N58)? \xnz.mem_r [779] : 
                        (N60)? \xnz.mem_r [812] : 
                        (N62)? \xnz.mem_r [845] : 
                        (N64)? \xnz.mem_r [878] : 
                        (N66)? \xnz.mem_r [911] : 
                        (N68)? \xnz.mem_r [944] : 
                        (N70)? \xnz.mem_r [977] : 
                        (N72)? \xnz.mem_r [1010] : 
                        (N74)? \xnz.mem_r [1043] : 1'b0;
  assign r_data_o[19] = (N43)? \xnz.mem_r [19] : 
                        (N45)? \xnz.mem_r [52] : 
                        (N47)? \xnz.mem_r [85] : 
                        (N49)? \xnz.mem_r [118] : 
                        (N51)? \xnz.mem_r [151] : 
                        (N53)? \xnz.mem_r [184] : 
                        (N55)? \xnz.mem_r [217] : 
                        (N57)? \xnz.mem_r [250] : 
                        (N59)? \xnz.mem_r [283] : 
                        (N61)? \xnz.mem_r [316] : 
                        (N63)? \xnz.mem_r [349] : 
                        (N65)? \xnz.mem_r [382] : 
                        (N67)? \xnz.mem_r [415] : 
                        (N69)? \xnz.mem_r [448] : 
                        (N71)? \xnz.mem_r [481] : 
                        (N73)? \xnz.mem_r [514] : 
                        (N44)? \xnz.mem_r [547] : 
                        (N46)? \xnz.mem_r [580] : 
                        (N48)? \xnz.mem_r [613] : 
                        (N50)? \xnz.mem_r [646] : 
                        (N52)? \xnz.mem_r [679] : 
                        (N54)? \xnz.mem_r [712] : 
                        (N56)? \xnz.mem_r [745] : 
                        (N58)? \xnz.mem_r [778] : 
                        (N60)? \xnz.mem_r [811] : 
                        (N62)? \xnz.mem_r [844] : 
                        (N64)? \xnz.mem_r [877] : 
                        (N66)? \xnz.mem_r [910] : 
                        (N68)? \xnz.mem_r [943] : 
                        (N70)? \xnz.mem_r [976] : 
                        (N72)? \xnz.mem_r [1009] : 
                        (N74)? \xnz.mem_r [1042] : 1'b0;
  assign r_data_o[18] = (N43)? \xnz.mem_r [18] : 
                        (N45)? \xnz.mem_r [51] : 
                        (N47)? \xnz.mem_r [84] : 
                        (N49)? \xnz.mem_r [117] : 
                        (N51)? \xnz.mem_r [150] : 
                        (N53)? \xnz.mem_r [183] : 
                        (N55)? \xnz.mem_r [216] : 
                        (N57)? \xnz.mem_r [249] : 
                        (N59)? \xnz.mem_r [282] : 
                        (N61)? \xnz.mem_r [315] : 
                        (N63)? \xnz.mem_r [348] : 
                        (N65)? \xnz.mem_r [381] : 
                        (N67)? \xnz.mem_r [414] : 
                        (N69)? \xnz.mem_r [447] : 
                        (N71)? \xnz.mem_r [480] : 
                        (N73)? \xnz.mem_r [513] : 
                        (N44)? \xnz.mem_r [546] : 
                        (N46)? \xnz.mem_r [579] : 
                        (N48)? \xnz.mem_r [612] : 
                        (N50)? \xnz.mem_r [645] : 
                        (N52)? \xnz.mem_r [678] : 
                        (N54)? \xnz.mem_r [711] : 
                        (N56)? \xnz.mem_r [744] : 
                        (N58)? \xnz.mem_r [777] : 
                        (N60)? \xnz.mem_r [810] : 
                        (N62)? \xnz.mem_r [843] : 
                        (N64)? \xnz.mem_r [876] : 
                        (N66)? \xnz.mem_r [909] : 
                        (N68)? \xnz.mem_r [942] : 
                        (N70)? \xnz.mem_r [975] : 
                        (N72)? \xnz.mem_r [1008] : 
                        (N74)? \xnz.mem_r [1041] : 1'b0;
  assign r_data_o[17] = (N43)? \xnz.mem_r [17] : 
                        (N45)? \xnz.mem_r [50] : 
                        (N47)? \xnz.mem_r [83] : 
                        (N49)? \xnz.mem_r [116] : 
                        (N51)? \xnz.mem_r [149] : 
                        (N53)? \xnz.mem_r [182] : 
                        (N55)? \xnz.mem_r [215] : 
                        (N57)? \xnz.mem_r [248] : 
                        (N59)? \xnz.mem_r [281] : 
                        (N61)? \xnz.mem_r [314] : 
                        (N63)? \xnz.mem_r [347] : 
                        (N65)? \xnz.mem_r [380] : 
                        (N67)? \xnz.mem_r [413] : 
                        (N69)? \xnz.mem_r [446] : 
                        (N71)? \xnz.mem_r [479] : 
                        (N73)? \xnz.mem_r [512] : 
                        (N44)? \xnz.mem_r [545] : 
                        (N46)? \xnz.mem_r [578] : 
                        (N48)? \xnz.mem_r [611] : 
                        (N50)? \xnz.mem_r [644] : 
                        (N52)? \xnz.mem_r [677] : 
                        (N54)? \xnz.mem_r [710] : 
                        (N56)? \xnz.mem_r [743] : 
                        (N58)? \xnz.mem_r [776] : 
                        (N60)? \xnz.mem_r [809] : 
                        (N62)? \xnz.mem_r [842] : 
                        (N64)? \xnz.mem_r [875] : 
                        (N66)? \xnz.mem_r [908] : 
                        (N68)? \xnz.mem_r [941] : 
                        (N70)? \xnz.mem_r [974] : 
                        (N72)? \xnz.mem_r [1007] : 
                        (N74)? \xnz.mem_r [1040] : 1'b0;
  assign r_data_o[16] = (N43)? \xnz.mem_r [16] : 
                        (N45)? \xnz.mem_r [49] : 
                        (N47)? \xnz.mem_r [82] : 
                        (N49)? \xnz.mem_r [115] : 
                        (N51)? \xnz.mem_r [148] : 
                        (N53)? \xnz.mem_r [181] : 
                        (N55)? \xnz.mem_r [214] : 
                        (N57)? \xnz.mem_r [247] : 
                        (N59)? \xnz.mem_r [280] : 
                        (N61)? \xnz.mem_r [313] : 
                        (N63)? \xnz.mem_r [346] : 
                        (N65)? \xnz.mem_r [379] : 
                        (N67)? \xnz.mem_r [412] : 
                        (N69)? \xnz.mem_r [445] : 
                        (N71)? \xnz.mem_r [478] : 
                        (N73)? \xnz.mem_r [511] : 
                        (N44)? \xnz.mem_r [544] : 
                        (N46)? \xnz.mem_r [577] : 
                        (N48)? \xnz.mem_r [610] : 
                        (N50)? \xnz.mem_r [643] : 
                        (N52)? \xnz.mem_r [676] : 
                        (N54)? \xnz.mem_r [709] : 
                        (N56)? \xnz.mem_r [742] : 
                        (N58)? \xnz.mem_r [775] : 
                        (N60)? \xnz.mem_r [808] : 
                        (N62)? \xnz.mem_r [841] : 
                        (N64)? \xnz.mem_r [874] : 
                        (N66)? \xnz.mem_r [907] : 
                        (N68)? \xnz.mem_r [940] : 
                        (N70)? \xnz.mem_r [973] : 
                        (N72)? \xnz.mem_r [1006] : 
                        (N74)? \xnz.mem_r [1039] : 1'b0;
  assign r_data_o[15] = (N43)? \xnz.mem_r [15] : 
                        (N45)? \xnz.mem_r [48] : 
                        (N47)? \xnz.mem_r [81] : 
                        (N49)? \xnz.mem_r [114] : 
                        (N51)? \xnz.mem_r [147] : 
                        (N53)? \xnz.mem_r [180] : 
                        (N55)? \xnz.mem_r [213] : 
                        (N57)? \xnz.mem_r [246] : 
                        (N59)? \xnz.mem_r [279] : 
                        (N61)? \xnz.mem_r [312] : 
                        (N63)? \xnz.mem_r [345] : 
                        (N65)? \xnz.mem_r [378] : 
                        (N67)? \xnz.mem_r [411] : 
                        (N69)? \xnz.mem_r [444] : 
                        (N71)? \xnz.mem_r [477] : 
                        (N73)? \xnz.mem_r [510] : 
                        (N44)? \xnz.mem_r [543] : 
                        (N46)? \xnz.mem_r [576] : 
                        (N48)? \xnz.mem_r [609] : 
                        (N50)? \xnz.mem_r [642] : 
                        (N52)? \xnz.mem_r [675] : 
                        (N54)? \xnz.mem_r [708] : 
                        (N56)? \xnz.mem_r [741] : 
                        (N58)? \xnz.mem_r [774] : 
                        (N60)? \xnz.mem_r [807] : 
                        (N62)? \xnz.mem_r [840] : 
                        (N64)? \xnz.mem_r [873] : 
                        (N66)? \xnz.mem_r [906] : 
                        (N68)? \xnz.mem_r [939] : 
                        (N70)? \xnz.mem_r [972] : 
                        (N72)? \xnz.mem_r [1005] : 
                        (N74)? \xnz.mem_r [1038] : 1'b0;
  assign r_data_o[14] = (N43)? \xnz.mem_r [14] : 
                        (N45)? \xnz.mem_r [47] : 
                        (N47)? \xnz.mem_r [80] : 
                        (N49)? \xnz.mem_r [113] : 
                        (N51)? \xnz.mem_r [146] : 
                        (N53)? \xnz.mem_r [179] : 
                        (N55)? \xnz.mem_r [212] : 
                        (N57)? \xnz.mem_r [245] : 
                        (N59)? \xnz.mem_r [278] : 
                        (N61)? \xnz.mem_r [311] : 
                        (N63)? \xnz.mem_r [344] : 
                        (N65)? \xnz.mem_r [377] : 
                        (N67)? \xnz.mem_r [410] : 
                        (N69)? \xnz.mem_r [443] : 
                        (N71)? \xnz.mem_r [476] : 
                        (N73)? \xnz.mem_r [509] : 
                        (N44)? \xnz.mem_r [542] : 
                        (N46)? \xnz.mem_r [575] : 
                        (N48)? \xnz.mem_r [608] : 
                        (N50)? \xnz.mem_r [641] : 
                        (N52)? \xnz.mem_r [674] : 
                        (N54)? \xnz.mem_r [707] : 
                        (N56)? \xnz.mem_r [740] : 
                        (N58)? \xnz.mem_r [773] : 
                        (N60)? \xnz.mem_r [806] : 
                        (N62)? \xnz.mem_r [839] : 
                        (N64)? \xnz.mem_r [872] : 
                        (N66)? \xnz.mem_r [905] : 
                        (N68)? \xnz.mem_r [938] : 
                        (N70)? \xnz.mem_r [971] : 
                        (N72)? \xnz.mem_r [1004] : 
                        (N74)? \xnz.mem_r [1037] : 1'b0;
  assign r_data_o[13] = (N43)? \xnz.mem_r [13] : 
                        (N45)? \xnz.mem_r [46] : 
                        (N47)? \xnz.mem_r [79] : 
                        (N49)? \xnz.mem_r [112] : 
                        (N51)? \xnz.mem_r [145] : 
                        (N53)? \xnz.mem_r [178] : 
                        (N55)? \xnz.mem_r [211] : 
                        (N57)? \xnz.mem_r [244] : 
                        (N59)? \xnz.mem_r [277] : 
                        (N61)? \xnz.mem_r [310] : 
                        (N63)? \xnz.mem_r [343] : 
                        (N65)? \xnz.mem_r [376] : 
                        (N67)? \xnz.mem_r [409] : 
                        (N69)? \xnz.mem_r [442] : 
                        (N71)? \xnz.mem_r [475] : 
                        (N73)? \xnz.mem_r [508] : 
                        (N44)? \xnz.mem_r [541] : 
                        (N46)? \xnz.mem_r [574] : 
                        (N48)? \xnz.mem_r [607] : 
                        (N50)? \xnz.mem_r [640] : 
                        (N52)? \xnz.mem_r [673] : 
                        (N54)? \xnz.mem_r [706] : 
                        (N56)? \xnz.mem_r [739] : 
                        (N58)? \xnz.mem_r [772] : 
                        (N60)? \xnz.mem_r [805] : 
                        (N62)? \xnz.mem_r [838] : 
                        (N64)? \xnz.mem_r [871] : 
                        (N66)? \xnz.mem_r [904] : 
                        (N68)? \xnz.mem_r [937] : 
                        (N70)? \xnz.mem_r [970] : 
                        (N72)? \xnz.mem_r [1003] : 
                        (N74)? \xnz.mem_r [1036] : 1'b0;
  assign r_data_o[12] = (N43)? \xnz.mem_r [12] : 
                        (N45)? \xnz.mem_r [45] : 
                        (N47)? \xnz.mem_r [78] : 
                        (N49)? \xnz.mem_r [111] : 
                        (N51)? \xnz.mem_r [144] : 
                        (N53)? \xnz.mem_r [177] : 
                        (N55)? \xnz.mem_r [210] : 
                        (N57)? \xnz.mem_r [243] : 
                        (N59)? \xnz.mem_r [276] : 
                        (N61)? \xnz.mem_r [309] : 
                        (N63)? \xnz.mem_r [342] : 
                        (N65)? \xnz.mem_r [375] : 
                        (N67)? \xnz.mem_r [408] : 
                        (N69)? \xnz.mem_r [441] : 
                        (N71)? \xnz.mem_r [474] : 
                        (N73)? \xnz.mem_r [507] : 
                        (N44)? \xnz.mem_r [540] : 
                        (N46)? \xnz.mem_r [573] : 
                        (N48)? \xnz.mem_r [606] : 
                        (N50)? \xnz.mem_r [639] : 
                        (N52)? \xnz.mem_r [672] : 
                        (N54)? \xnz.mem_r [705] : 
                        (N56)? \xnz.mem_r [738] : 
                        (N58)? \xnz.mem_r [771] : 
                        (N60)? \xnz.mem_r [804] : 
                        (N62)? \xnz.mem_r [837] : 
                        (N64)? \xnz.mem_r [870] : 
                        (N66)? \xnz.mem_r [903] : 
                        (N68)? \xnz.mem_r [936] : 
                        (N70)? \xnz.mem_r [969] : 
                        (N72)? \xnz.mem_r [1002] : 
                        (N74)? \xnz.mem_r [1035] : 1'b0;
  assign r_data_o[11] = (N43)? \xnz.mem_r [11] : 
                        (N45)? \xnz.mem_r [44] : 
                        (N47)? \xnz.mem_r [77] : 
                        (N49)? \xnz.mem_r [110] : 
                        (N51)? \xnz.mem_r [143] : 
                        (N53)? \xnz.mem_r [176] : 
                        (N55)? \xnz.mem_r [209] : 
                        (N57)? \xnz.mem_r [242] : 
                        (N59)? \xnz.mem_r [275] : 
                        (N61)? \xnz.mem_r [308] : 
                        (N63)? \xnz.mem_r [341] : 
                        (N65)? \xnz.mem_r [374] : 
                        (N67)? \xnz.mem_r [407] : 
                        (N69)? \xnz.mem_r [440] : 
                        (N71)? \xnz.mem_r [473] : 
                        (N73)? \xnz.mem_r [506] : 
                        (N44)? \xnz.mem_r [539] : 
                        (N46)? \xnz.mem_r [572] : 
                        (N48)? \xnz.mem_r [605] : 
                        (N50)? \xnz.mem_r [638] : 
                        (N52)? \xnz.mem_r [671] : 
                        (N54)? \xnz.mem_r [704] : 
                        (N56)? \xnz.mem_r [737] : 
                        (N58)? \xnz.mem_r [770] : 
                        (N60)? \xnz.mem_r [803] : 
                        (N62)? \xnz.mem_r [836] : 
                        (N64)? \xnz.mem_r [869] : 
                        (N66)? \xnz.mem_r [902] : 
                        (N68)? \xnz.mem_r [935] : 
                        (N70)? \xnz.mem_r [968] : 
                        (N72)? \xnz.mem_r [1001] : 
                        (N74)? \xnz.mem_r [1034] : 1'b0;
  assign r_data_o[10] = (N43)? \xnz.mem_r [10] : 
                        (N45)? \xnz.mem_r [43] : 
                        (N47)? \xnz.mem_r [76] : 
                        (N49)? \xnz.mem_r [109] : 
                        (N51)? \xnz.mem_r [142] : 
                        (N53)? \xnz.mem_r [175] : 
                        (N55)? \xnz.mem_r [208] : 
                        (N57)? \xnz.mem_r [241] : 
                        (N59)? \xnz.mem_r [274] : 
                        (N61)? \xnz.mem_r [307] : 
                        (N63)? \xnz.mem_r [340] : 
                        (N65)? \xnz.mem_r [373] : 
                        (N67)? \xnz.mem_r [406] : 
                        (N69)? \xnz.mem_r [439] : 
                        (N71)? \xnz.mem_r [472] : 
                        (N73)? \xnz.mem_r [505] : 
                        (N44)? \xnz.mem_r [538] : 
                        (N46)? \xnz.mem_r [571] : 
                        (N48)? \xnz.mem_r [604] : 
                        (N50)? \xnz.mem_r [637] : 
                        (N52)? \xnz.mem_r [670] : 
                        (N54)? \xnz.mem_r [703] : 
                        (N56)? \xnz.mem_r [736] : 
                        (N58)? \xnz.mem_r [769] : 
                        (N60)? \xnz.mem_r [802] : 
                        (N62)? \xnz.mem_r [835] : 
                        (N64)? \xnz.mem_r [868] : 
                        (N66)? \xnz.mem_r [901] : 
                        (N68)? \xnz.mem_r [934] : 
                        (N70)? \xnz.mem_r [967] : 
                        (N72)? \xnz.mem_r [1000] : 
                        (N74)? \xnz.mem_r [1033] : 1'b0;
  assign r_data_o[9] = (N43)? \xnz.mem_r [9] : 
                       (N45)? \xnz.mem_r [42] : 
                       (N47)? \xnz.mem_r [75] : 
                       (N49)? \xnz.mem_r [108] : 
                       (N51)? \xnz.mem_r [141] : 
                       (N53)? \xnz.mem_r [174] : 
                       (N55)? \xnz.mem_r [207] : 
                       (N57)? \xnz.mem_r [240] : 
                       (N59)? \xnz.mem_r [273] : 
                       (N61)? \xnz.mem_r [306] : 
                       (N63)? \xnz.mem_r [339] : 
                       (N65)? \xnz.mem_r [372] : 
                       (N67)? \xnz.mem_r [405] : 
                       (N69)? \xnz.mem_r [438] : 
                       (N71)? \xnz.mem_r [471] : 
                       (N73)? \xnz.mem_r [504] : 
                       (N44)? \xnz.mem_r [537] : 
                       (N46)? \xnz.mem_r [570] : 
                       (N48)? \xnz.mem_r [603] : 
                       (N50)? \xnz.mem_r [636] : 
                       (N52)? \xnz.mem_r [669] : 
                       (N54)? \xnz.mem_r [702] : 
                       (N56)? \xnz.mem_r [735] : 
                       (N58)? \xnz.mem_r [768] : 
                       (N60)? \xnz.mem_r [801] : 
                       (N62)? \xnz.mem_r [834] : 
                       (N64)? \xnz.mem_r [867] : 
                       (N66)? \xnz.mem_r [900] : 
                       (N68)? \xnz.mem_r [933] : 
                       (N70)? \xnz.mem_r [966] : 
                       (N72)? \xnz.mem_r [999] : 
                       (N74)? \xnz.mem_r [1032] : 1'b0;
  assign r_data_o[8] = (N43)? \xnz.mem_r [8] : 
                       (N45)? \xnz.mem_r [41] : 
                       (N47)? \xnz.mem_r [74] : 
                       (N49)? \xnz.mem_r [107] : 
                       (N51)? \xnz.mem_r [140] : 
                       (N53)? \xnz.mem_r [173] : 
                       (N55)? \xnz.mem_r [206] : 
                       (N57)? \xnz.mem_r [239] : 
                       (N59)? \xnz.mem_r [272] : 
                       (N61)? \xnz.mem_r [305] : 
                       (N63)? \xnz.mem_r [338] : 
                       (N65)? \xnz.mem_r [371] : 
                       (N67)? \xnz.mem_r [404] : 
                       (N69)? \xnz.mem_r [437] : 
                       (N71)? \xnz.mem_r [470] : 
                       (N73)? \xnz.mem_r [503] : 
                       (N44)? \xnz.mem_r [536] : 
                       (N46)? \xnz.mem_r [569] : 
                       (N48)? \xnz.mem_r [602] : 
                       (N50)? \xnz.mem_r [635] : 
                       (N52)? \xnz.mem_r [668] : 
                       (N54)? \xnz.mem_r [701] : 
                       (N56)? \xnz.mem_r [734] : 
                       (N58)? \xnz.mem_r [767] : 
                       (N60)? \xnz.mem_r [800] : 
                       (N62)? \xnz.mem_r [833] : 
                       (N64)? \xnz.mem_r [866] : 
                       (N66)? \xnz.mem_r [899] : 
                       (N68)? \xnz.mem_r [932] : 
                       (N70)? \xnz.mem_r [965] : 
                       (N72)? \xnz.mem_r [998] : 
                       (N74)? \xnz.mem_r [1031] : 1'b0;
  assign r_data_o[7] = (N43)? \xnz.mem_r [7] : 
                       (N45)? \xnz.mem_r [40] : 
                       (N47)? \xnz.mem_r [73] : 
                       (N49)? \xnz.mem_r [106] : 
                       (N51)? \xnz.mem_r [139] : 
                       (N53)? \xnz.mem_r [172] : 
                       (N55)? \xnz.mem_r [205] : 
                       (N57)? \xnz.mem_r [238] : 
                       (N59)? \xnz.mem_r [271] : 
                       (N61)? \xnz.mem_r [304] : 
                       (N63)? \xnz.mem_r [337] : 
                       (N65)? \xnz.mem_r [370] : 
                       (N67)? \xnz.mem_r [403] : 
                       (N69)? \xnz.mem_r [436] : 
                       (N71)? \xnz.mem_r [469] : 
                       (N73)? \xnz.mem_r [502] : 
                       (N44)? \xnz.mem_r [535] : 
                       (N46)? \xnz.mem_r [568] : 
                       (N48)? \xnz.mem_r [601] : 
                       (N50)? \xnz.mem_r [634] : 
                       (N52)? \xnz.mem_r [667] : 
                       (N54)? \xnz.mem_r [700] : 
                       (N56)? \xnz.mem_r [733] : 
                       (N58)? \xnz.mem_r [766] : 
                       (N60)? \xnz.mem_r [799] : 
                       (N62)? \xnz.mem_r [832] : 
                       (N64)? \xnz.mem_r [865] : 
                       (N66)? \xnz.mem_r [898] : 
                       (N68)? \xnz.mem_r [931] : 
                       (N70)? \xnz.mem_r [964] : 
                       (N72)? \xnz.mem_r [997] : 
                       (N74)? \xnz.mem_r [1030] : 1'b0;
  assign r_data_o[6] = (N43)? \xnz.mem_r [6] : 
                       (N45)? \xnz.mem_r [39] : 
                       (N47)? \xnz.mem_r [72] : 
                       (N49)? \xnz.mem_r [105] : 
                       (N51)? \xnz.mem_r [138] : 
                       (N53)? \xnz.mem_r [171] : 
                       (N55)? \xnz.mem_r [204] : 
                       (N57)? \xnz.mem_r [237] : 
                       (N59)? \xnz.mem_r [270] : 
                       (N61)? \xnz.mem_r [303] : 
                       (N63)? \xnz.mem_r [336] : 
                       (N65)? \xnz.mem_r [369] : 
                       (N67)? \xnz.mem_r [402] : 
                       (N69)? \xnz.mem_r [435] : 
                       (N71)? \xnz.mem_r [468] : 
                       (N73)? \xnz.mem_r [501] : 
                       (N44)? \xnz.mem_r [534] : 
                       (N46)? \xnz.mem_r [567] : 
                       (N48)? \xnz.mem_r [600] : 
                       (N50)? \xnz.mem_r [633] : 
                       (N52)? \xnz.mem_r [666] : 
                       (N54)? \xnz.mem_r [699] : 
                       (N56)? \xnz.mem_r [732] : 
                       (N58)? \xnz.mem_r [765] : 
                       (N60)? \xnz.mem_r [798] : 
                       (N62)? \xnz.mem_r [831] : 
                       (N64)? \xnz.mem_r [864] : 
                       (N66)? \xnz.mem_r [897] : 
                       (N68)? \xnz.mem_r [930] : 
                       (N70)? \xnz.mem_r [963] : 
                       (N72)? \xnz.mem_r [996] : 
                       (N74)? \xnz.mem_r [1029] : 1'b0;
  assign r_data_o[5] = (N43)? \xnz.mem_r [5] : 
                       (N45)? \xnz.mem_r [38] : 
                       (N47)? \xnz.mem_r [71] : 
                       (N49)? \xnz.mem_r [104] : 
                       (N51)? \xnz.mem_r [137] : 
                       (N53)? \xnz.mem_r [170] : 
                       (N55)? \xnz.mem_r [203] : 
                       (N57)? \xnz.mem_r [236] : 
                       (N59)? \xnz.mem_r [269] : 
                       (N61)? \xnz.mem_r [302] : 
                       (N63)? \xnz.mem_r [335] : 
                       (N65)? \xnz.mem_r [368] : 
                       (N67)? \xnz.mem_r [401] : 
                       (N69)? \xnz.mem_r [434] : 
                       (N71)? \xnz.mem_r [467] : 
                       (N73)? \xnz.mem_r [500] : 
                       (N44)? \xnz.mem_r [533] : 
                       (N46)? \xnz.mem_r [566] : 
                       (N48)? \xnz.mem_r [599] : 
                       (N50)? \xnz.mem_r [632] : 
                       (N52)? \xnz.mem_r [665] : 
                       (N54)? \xnz.mem_r [698] : 
                       (N56)? \xnz.mem_r [731] : 
                       (N58)? \xnz.mem_r [764] : 
                       (N60)? \xnz.mem_r [797] : 
                       (N62)? \xnz.mem_r [830] : 
                       (N64)? \xnz.mem_r [863] : 
                       (N66)? \xnz.mem_r [896] : 
                       (N68)? \xnz.mem_r [929] : 
                       (N70)? \xnz.mem_r [962] : 
                       (N72)? \xnz.mem_r [995] : 
                       (N74)? \xnz.mem_r [1028] : 1'b0;
  assign r_data_o[4] = (N43)? \xnz.mem_r [4] : 
                       (N45)? \xnz.mem_r [37] : 
                       (N47)? \xnz.mem_r [70] : 
                       (N49)? \xnz.mem_r [103] : 
                       (N51)? \xnz.mem_r [136] : 
                       (N53)? \xnz.mem_r [169] : 
                       (N55)? \xnz.mem_r [202] : 
                       (N57)? \xnz.mem_r [235] : 
                       (N59)? \xnz.mem_r [268] : 
                       (N61)? \xnz.mem_r [301] : 
                       (N63)? \xnz.mem_r [334] : 
                       (N65)? \xnz.mem_r [367] : 
                       (N67)? \xnz.mem_r [400] : 
                       (N69)? \xnz.mem_r [433] : 
                       (N71)? \xnz.mem_r [466] : 
                       (N73)? \xnz.mem_r [499] : 
                       (N44)? \xnz.mem_r [532] : 
                       (N46)? \xnz.mem_r [565] : 
                       (N48)? \xnz.mem_r [598] : 
                       (N50)? \xnz.mem_r [631] : 
                       (N52)? \xnz.mem_r [664] : 
                       (N54)? \xnz.mem_r [697] : 
                       (N56)? \xnz.mem_r [730] : 
                       (N58)? \xnz.mem_r [763] : 
                       (N60)? \xnz.mem_r [796] : 
                       (N62)? \xnz.mem_r [829] : 
                       (N64)? \xnz.mem_r [862] : 
                       (N66)? \xnz.mem_r [895] : 
                       (N68)? \xnz.mem_r [928] : 
                       (N70)? \xnz.mem_r [961] : 
                       (N72)? \xnz.mem_r [994] : 
                       (N74)? \xnz.mem_r [1027] : 1'b0;
  assign r_data_o[3] = (N43)? \xnz.mem_r [3] : 
                       (N45)? \xnz.mem_r [36] : 
                       (N47)? \xnz.mem_r [69] : 
                       (N49)? \xnz.mem_r [102] : 
                       (N51)? \xnz.mem_r [135] : 
                       (N53)? \xnz.mem_r [168] : 
                       (N55)? \xnz.mem_r [201] : 
                       (N57)? \xnz.mem_r [234] : 
                       (N59)? \xnz.mem_r [267] : 
                       (N61)? \xnz.mem_r [300] : 
                       (N63)? \xnz.mem_r [333] : 
                       (N65)? \xnz.mem_r [366] : 
                       (N67)? \xnz.mem_r [399] : 
                       (N69)? \xnz.mem_r [432] : 
                       (N71)? \xnz.mem_r [465] : 
                       (N73)? \xnz.mem_r [498] : 
                       (N44)? \xnz.mem_r [531] : 
                       (N46)? \xnz.mem_r [564] : 
                       (N48)? \xnz.mem_r [597] : 
                       (N50)? \xnz.mem_r [630] : 
                       (N52)? \xnz.mem_r [663] : 
                       (N54)? \xnz.mem_r [696] : 
                       (N56)? \xnz.mem_r [729] : 
                       (N58)? \xnz.mem_r [762] : 
                       (N60)? \xnz.mem_r [795] : 
                       (N62)? \xnz.mem_r [828] : 
                       (N64)? \xnz.mem_r [861] : 
                       (N66)? \xnz.mem_r [894] : 
                       (N68)? \xnz.mem_r [927] : 
                       (N70)? \xnz.mem_r [960] : 
                       (N72)? \xnz.mem_r [993] : 
                       (N74)? \xnz.mem_r [1026] : 1'b0;
  assign r_data_o[2] = (N43)? \xnz.mem_r [2] : 
                       (N45)? \xnz.mem_r [35] : 
                       (N47)? \xnz.mem_r [68] : 
                       (N49)? \xnz.mem_r [101] : 
                       (N51)? \xnz.mem_r [134] : 
                       (N53)? \xnz.mem_r [167] : 
                       (N55)? \xnz.mem_r [200] : 
                       (N57)? \xnz.mem_r [233] : 
                       (N59)? \xnz.mem_r [266] : 
                       (N61)? \xnz.mem_r [299] : 
                       (N63)? \xnz.mem_r [332] : 
                       (N65)? \xnz.mem_r [365] : 
                       (N67)? \xnz.mem_r [398] : 
                       (N69)? \xnz.mem_r [431] : 
                       (N71)? \xnz.mem_r [464] : 
                       (N73)? \xnz.mem_r [497] : 
                       (N44)? \xnz.mem_r [530] : 
                       (N46)? \xnz.mem_r [563] : 
                       (N48)? \xnz.mem_r [596] : 
                       (N50)? \xnz.mem_r [629] : 
                       (N52)? \xnz.mem_r [662] : 
                       (N54)? \xnz.mem_r [695] : 
                       (N56)? \xnz.mem_r [728] : 
                       (N58)? \xnz.mem_r [761] : 
                       (N60)? \xnz.mem_r [794] : 
                       (N62)? \xnz.mem_r [827] : 
                       (N64)? \xnz.mem_r [860] : 
                       (N66)? \xnz.mem_r [893] : 
                       (N68)? \xnz.mem_r [926] : 
                       (N70)? \xnz.mem_r [959] : 
                       (N72)? \xnz.mem_r [992] : 
                       (N74)? \xnz.mem_r [1025] : 1'b0;
  assign r_data_o[1] = (N43)? \xnz.mem_r [1] : 
                       (N45)? \xnz.mem_r [34] : 
                       (N47)? \xnz.mem_r [67] : 
                       (N49)? \xnz.mem_r [100] : 
                       (N51)? \xnz.mem_r [133] : 
                       (N53)? \xnz.mem_r [166] : 
                       (N55)? \xnz.mem_r [199] : 
                       (N57)? \xnz.mem_r [232] : 
                       (N59)? \xnz.mem_r [265] : 
                       (N61)? \xnz.mem_r [298] : 
                       (N63)? \xnz.mem_r [331] : 
                       (N65)? \xnz.mem_r [364] : 
                       (N67)? \xnz.mem_r [397] : 
                       (N69)? \xnz.mem_r [430] : 
                       (N71)? \xnz.mem_r [463] : 
                       (N73)? \xnz.mem_r [496] : 
                       (N44)? \xnz.mem_r [529] : 
                       (N46)? \xnz.mem_r [562] : 
                       (N48)? \xnz.mem_r [595] : 
                       (N50)? \xnz.mem_r [628] : 
                       (N52)? \xnz.mem_r [661] : 
                       (N54)? \xnz.mem_r [694] : 
                       (N56)? \xnz.mem_r [727] : 
                       (N58)? \xnz.mem_r [760] : 
                       (N60)? \xnz.mem_r [793] : 
                       (N62)? \xnz.mem_r [826] : 
                       (N64)? \xnz.mem_r [859] : 
                       (N66)? \xnz.mem_r [892] : 
                       (N68)? \xnz.mem_r [925] : 
                       (N70)? \xnz.mem_r [958] : 
                       (N72)? \xnz.mem_r [991] : 
                       (N74)? \xnz.mem_r [1024] : 1'b0;
  assign r_data_o[0] = (N43)? \xnz.mem_r [0] : 
                       (N45)? \xnz.mem_r [33] : 
                       (N47)? \xnz.mem_r [66] : 
                       (N49)? \xnz.mem_r [99] : 
                       (N51)? \xnz.mem_r [132] : 
                       (N53)? \xnz.mem_r [165] : 
                       (N55)? \xnz.mem_r [198] : 
                       (N57)? \xnz.mem_r [231] : 
                       (N59)? \xnz.mem_r [264] : 
                       (N61)? \xnz.mem_r [297] : 
                       (N63)? \xnz.mem_r [330] : 
                       (N65)? \xnz.mem_r [363] : 
                       (N67)? \xnz.mem_r [396] : 
                       (N69)? \xnz.mem_r [429] : 
                       (N71)? \xnz.mem_r [462] : 
                       (N73)? \xnz.mem_r [495] : 
                       (N44)? \xnz.mem_r [528] : 
                       (N46)? \xnz.mem_r [561] : 
                       (N48)? \xnz.mem_r [594] : 
                       (N50)? \xnz.mem_r [627] : 
                       (N52)? \xnz.mem_r [660] : 
                       (N54)? \xnz.mem_r [693] : 
                       (N56)? \xnz.mem_r [726] : 
                       (N58)? \xnz.mem_r [759] : 
                       (N60)? \xnz.mem_r [792] : 
                       (N62)? \xnz.mem_r [825] : 
                       (N64)? \xnz.mem_r [858] : 
                       (N66)? \xnz.mem_r [891] : 
                       (N68)? \xnz.mem_r [924] : 
                       (N70)? \xnz.mem_r [957] : 
                       (N72)? \xnz.mem_r [990] : 
                       (N74)? \xnz.mem_r [1023] : 1'b0;
  assign r_data_o[65] = (N108)? \xnz.mem_r [32] : 
                        (N110)? \xnz.mem_r [65] : 
                        (N112)? \xnz.mem_r [98] : 
                        (N114)? \xnz.mem_r [131] : 
                        (N116)? \xnz.mem_r [164] : 
                        (N118)? \xnz.mem_r [197] : 
                        (N120)? \xnz.mem_r [230] : 
                        (N122)? \xnz.mem_r [263] : 
                        (N124)? \xnz.mem_r [296] : 
                        (N126)? \xnz.mem_r [329] : 
                        (N128)? \xnz.mem_r [362] : 
                        (N130)? \xnz.mem_r [395] : 
                        (N132)? \xnz.mem_r [428] : 
                        (N134)? \xnz.mem_r [461] : 
                        (N136)? \xnz.mem_r [494] : 
                        (N138)? \xnz.mem_r [527] : 
                        (N109)? \xnz.mem_r [560] : 
                        (N111)? \xnz.mem_r [593] : 
                        (N113)? \xnz.mem_r [626] : 
                        (N115)? \xnz.mem_r [659] : 
                        (N117)? \xnz.mem_r [692] : 
                        (N119)? \xnz.mem_r [725] : 
                        (N121)? \xnz.mem_r [758] : 
                        (N123)? \xnz.mem_r [791] : 
                        (N125)? \xnz.mem_r [824] : 
                        (N127)? \xnz.mem_r [857] : 
                        (N129)? \xnz.mem_r [890] : 
                        (N131)? \xnz.mem_r [923] : 
                        (N133)? \xnz.mem_r [956] : 
                        (N135)? \xnz.mem_r [989] : 
                        (N137)? \xnz.mem_r [1022] : 
                        (N139)? \xnz.mem_r [1055] : 1'b0;
  assign r_data_o[64] = (N108)? \xnz.mem_r [31] : 
                        (N110)? \xnz.mem_r [64] : 
                        (N112)? \xnz.mem_r [97] : 
                        (N114)? \xnz.mem_r [130] : 
                        (N116)? \xnz.mem_r [163] : 
                        (N118)? \xnz.mem_r [196] : 
                        (N120)? \xnz.mem_r [229] : 
                        (N122)? \xnz.mem_r [262] : 
                        (N124)? \xnz.mem_r [295] : 
                        (N126)? \xnz.mem_r [328] : 
                        (N128)? \xnz.mem_r [361] : 
                        (N130)? \xnz.mem_r [394] : 
                        (N132)? \xnz.mem_r [427] : 
                        (N134)? \xnz.mem_r [460] : 
                        (N136)? \xnz.mem_r [493] : 
                        (N138)? \xnz.mem_r [526] : 
                        (N109)? \xnz.mem_r [559] : 
                        (N111)? \xnz.mem_r [592] : 
                        (N113)? \xnz.mem_r [625] : 
                        (N115)? \xnz.mem_r [658] : 
                        (N117)? \xnz.mem_r [691] : 
                        (N119)? \xnz.mem_r [724] : 
                        (N121)? \xnz.mem_r [757] : 
                        (N123)? \xnz.mem_r [790] : 
                        (N125)? \xnz.mem_r [823] : 
                        (N127)? \xnz.mem_r [856] : 
                        (N129)? \xnz.mem_r [889] : 
                        (N131)? \xnz.mem_r [922] : 
                        (N133)? \xnz.mem_r [955] : 
                        (N135)? \xnz.mem_r [988] : 
                        (N137)? \xnz.mem_r [1021] : 
                        (N139)? \xnz.mem_r [1054] : 1'b0;
  assign r_data_o[63] = (N108)? \xnz.mem_r [30] : 
                        (N110)? \xnz.mem_r [63] : 
                        (N112)? \xnz.mem_r [96] : 
                        (N114)? \xnz.mem_r [129] : 
                        (N116)? \xnz.mem_r [162] : 
                        (N118)? \xnz.mem_r [195] : 
                        (N120)? \xnz.mem_r [228] : 
                        (N122)? \xnz.mem_r [261] : 
                        (N124)? \xnz.mem_r [294] : 
                        (N126)? \xnz.mem_r [327] : 
                        (N128)? \xnz.mem_r [360] : 
                        (N130)? \xnz.mem_r [393] : 
                        (N132)? \xnz.mem_r [426] : 
                        (N134)? \xnz.mem_r [459] : 
                        (N136)? \xnz.mem_r [492] : 
                        (N138)? \xnz.mem_r [525] : 
                        (N109)? \xnz.mem_r [558] : 
                        (N111)? \xnz.mem_r [591] : 
                        (N113)? \xnz.mem_r [624] : 
                        (N115)? \xnz.mem_r [657] : 
                        (N117)? \xnz.mem_r [690] : 
                        (N119)? \xnz.mem_r [723] : 
                        (N121)? \xnz.mem_r [756] : 
                        (N123)? \xnz.mem_r [789] : 
                        (N125)? \xnz.mem_r [822] : 
                        (N127)? \xnz.mem_r [855] : 
                        (N129)? \xnz.mem_r [888] : 
                        (N131)? \xnz.mem_r [921] : 
                        (N133)? \xnz.mem_r [954] : 
                        (N135)? \xnz.mem_r [987] : 
                        (N137)? \xnz.mem_r [1020] : 
                        (N139)? \xnz.mem_r [1053] : 1'b0;
  assign r_data_o[62] = (N108)? \xnz.mem_r [29] : 
                        (N110)? \xnz.mem_r [62] : 
                        (N112)? \xnz.mem_r [95] : 
                        (N114)? \xnz.mem_r [128] : 
                        (N116)? \xnz.mem_r [161] : 
                        (N118)? \xnz.mem_r [194] : 
                        (N120)? \xnz.mem_r [227] : 
                        (N122)? \xnz.mem_r [260] : 
                        (N124)? \xnz.mem_r [293] : 
                        (N126)? \xnz.mem_r [326] : 
                        (N128)? \xnz.mem_r [359] : 
                        (N130)? \xnz.mem_r [392] : 
                        (N132)? \xnz.mem_r [425] : 
                        (N134)? \xnz.mem_r [458] : 
                        (N136)? \xnz.mem_r [491] : 
                        (N138)? \xnz.mem_r [524] : 
                        (N109)? \xnz.mem_r [557] : 
                        (N111)? \xnz.mem_r [590] : 
                        (N113)? \xnz.mem_r [623] : 
                        (N115)? \xnz.mem_r [656] : 
                        (N117)? \xnz.mem_r [689] : 
                        (N119)? \xnz.mem_r [722] : 
                        (N121)? \xnz.mem_r [755] : 
                        (N123)? \xnz.mem_r [788] : 
                        (N125)? \xnz.mem_r [821] : 
                        (N127)? \xnz.mem_r [854] : 
                        (N129)? \xnz.mem_r [887] : 
                        (N131)? \xnz.mem_r [920] : 
                        (N133)? \xnz.mem_r [953] : 
                        (N135)? \xnz.mem_r [986] : 
                        (N137)? \xnz.mem_r [1019] : 
                        (N139)? \xnz.mem_r [1052] : 1'b0;
  assign r_data_o[61] = (N108)? \xnz.mem_r [28] : 
                        (N110)? \xnz.mem_r [61] : 
                        (N112)? \xnz.mem_r [94] : 
                        (N114)? \xnz.mem_r [127] : 
                        (N116)? \xnz.mem_r [160] : 
                        (N118)? \xnz.mem_r [193] : 
                        (N120)? \xnz.mem_r [226] : 
                        (N122)? \xnz.mem_r [259] : 
                        (N124)? \xnz.mem_r [292] : 
                        (N126)? \xnz.mem_r [325] : 
                        (N128)? \xnz.mem_r [358] : 
                        (N130)? \xnz.mem_r [391] : 
                        (N132)? \xnz.mem_r [424] : 
                        (N134)? \xnz.mem_r [457] : 
                        (N136)? \xnz.mem_r [490] : 
                        (N138)? \xnz.mem_r [523] : 
                        (N109)? \xnz.mem_r [556] : 
                        (N111)? \xnz.mem_r [589] : 
                        (N113)? \xnz.mem_r [622] : 
                        (N115)? \xnz.mem_r [655] : 
                        (N117)? \xnz.mem_r [688] : 
                        (N119)? \xnz.mem_r [721] : 
                        (N121)? \xnz.mem_r [754] : 
                        (N123)? \xnz.mem_r [787] : 
                        (N125)? \xnz.mem_r [820] : 
                        (N127)? \xnz.mem_r [853] : 
                        (N129)? \xnz.mem_r [886] : 
                        (N131)? \xnz.mem_r [919] : 
                        (N133)? \xnz.mem_r [952] : 
                        (N135)? \xnz.mem_r [985] : 
                        (N137)? \xnz.mem_r [1018] : 
                        (N139)? \xnz.mem_r [1051] : 1'b0;
  assign r_data_o[60] = (N108)? \xnz.mem_r [27] : 
                        (N110)? \xnz.mem_r [60] : 
                        (N112)? \xnz.mem_r [93] : 
                        (N114)? \xnz.mem_r [126] : 
                        (N116)? \xnz.mem_r [159] : 
                        (N118)? \xnz.mem_r [192] : 
                        (N120)? \xnz.mem_r [225] : 
                        (N122)? \xnz.mem_r [258] : 
                        (N124)? \xnz.mem_r [291] : 
                        (N126)? \xnz.mem_r [324] : 
                        (N128)? \xnz.mem_r [357] : 
                        (N130)? \xnz.mem_r [390] : 
                        (N132)? \xnz.mem_r [423] : 
                        (N134)? \xnz.mem_r [456] : 
                        (N136)? \xnz.mem_r [489] : 
                        (N138)? \xnz.mem_r [522] : 
                        (N109)? \xnz.mem_r [555] : 
                        (N111)? \xnz.mem_r [588] : 
                        (N113)? \xnz.mem_r [621] : 
                        (N115)? \xnz.mem_r [654] : 
                        (N117)? \xnz.mem_r [687] : 
                        (N119)? \xnz.mem_r [720] : 
                        (N121)? \xnz.mem_r [753] : 
                        (N123)? \xnz.mem_r [786] : 
                        (N125)? \xnz.mem_r [819] : 
                        (N127)? \xnz.mem_r [852] : 
                        (N129)? \xnz.mem_r [885] : 
                        (N131)? \xnz.mem_r [918] : 
                        (N133)? \xnz.mem_r [951] : 
                        (N135)? \xnz.mem_r [984] : 
                        (N137)? \xnz.mem_r [1017] : 
                        (N139)? \xnz.mem_r [1050] : 1'b0;
  assign r_data_o[59] = (N108)? \xnz.mem_r [26] : 
                        (N110)? \xnz.mem_r [59] : 
                        (N112)? \xnz.mem_r [92] : 
                        (N114)? \xnz.mem_r [125] : 
                        (N116)? \xnz.mem_r [158] : 
                        (N118)? \xnz.mem_r [191] : 
                        (N120)? \xnz.mem_r [224] : 
                        (N122)? \xnz.mem_r [257] : 
                        (N124)? \xnz.mem_r [290] : 
                        (N126)? \xnz.mem_r [323] : 
                        (N128)? \xnz.mem_r [356] : 
                        (N130)? \xnz.mem_r [389] : 
                        (N132)? \xnz.mem_r [422] : 
                        (N134)? \xnz.mem_r [455] : 
                        (N136)? \xnz.mem_r [488] : 
                        (N138)? \xnz.mem_r [521] : 
                        (N109)? \xnz.mem_r [554] : 
                        (N111)? \xnz.mem_r [587] : 
                        (N113)? \xnz.mem_r [620] : 
                        (N115)? \xnz.mem_r [653] : 
                        (N117)? \xnz.mem_r [686] : 
                        (N119)? \xnz.mem_r [719] : 
                        (N121)? \xnz.mem_r [752] : 
                        (N123)? \xnz.mem_r [785] : 
                        (N125)? \xnz.mem_r [818] : 
                        (N127)? \xnz.mem_r [851] : 
                        (N129)? \xnz.mem_r [884] : 
                        (N131)? \xnz.mem_r [917] : 
                        (N133)? \xnz.mem_r [950] : 
                        (N135)? \xnz.mem_r [983] : 
                        (N137)? \xnz.mem_r [1016] : 
                        (N139)? \xnz.mem_r [1049] : 1'b0;
  assign r_data_o[58] = (N108)? \xnz.mem_r [25] : 
                        (N110)? \xnz.mem_r [58] : 
                        (N112)? \xnz.mem_r [91] : 
                        (N114)? \xnz.mem_r [124] : 
                        (N116)? \xnz.mem_r [157] : 
                        (N118)? \xnz.mem_r [190] : 
                        (N120)? \xnz.mem_r [223] : 
                        (N122)? \xnz.mem_r [256] : 
                        (N124)? \xnz.mem_r [289] : 
                        (N126)? \xnz.mem_r [322] : 
                        (N128)? \xnz.mem_r [355] : 
                        (N130)? \xnz.mem_r [388] : 
                        (N132)? \xnz.mem_r [421] : 
                        (N134)? \xnz.mem_r [454] : 
                        (N136)? \xnz.mem_r [487] : 
                        (N138)? \xnz.mem_r [520] : 
                        (N109)? \xnz.mem_r [553] : 
                        (N111)? \xnz.mem_r [586] : 
                        (N113)? \xnz.mem_r [619] : 
                        (N115)? \xnz.mem_r [652] : 
                        (N117)? \xnz.mem_r [685] : 
                        (N119)? \xnz.mem_r [718] : 
                        (N121)? \xnz.mem_r [751] : 
                        (N123)? \xnz.mem_r [784] : 
                        (N125)? \xnz.mem_r [817] : 
                        (N127)? \xnz.mem_r [850] : 
                        (N129)? \xnz.mem_r [883] : 
                        (N131)? \xnz.mem_r [916] : 
                        (N133)? \xnz.mem_r [949] : 
                        (N135)? \xnz.mem_r [982] : 
                        (N137)? \xnz.mem_r [1015] : 
                        (N139)? \xnz.mem_r [1048] : 1'b0;
  assign r_data_o[57] = (N108)? \xnz.mem_r [24] : 
                        (N110)? \xnz.mem_r [57] : 
                        (N112)? \xnz.mem_r [90] : 
                        (N114)? \xnz.mem_r [123] : 
                        (N116)? \xnz.mem_r [156] : 
                        (N118)? \xnz.mem_r [189] : 
                        (N120)? \xnz.mem_r [222] : 
                        (N122)? \xnz.mem_r [255] : 
                        (N124)? \xnz.mem_r [288] : 
                        (N126)? \xnz.mem_r [321] : 
                        (N128)? \xnz.mem_r [354] : 
                        (N130)? \xnz.mem_r [387] : 
                        (N132)? \xnz.mem_r [420] : 
                        (N134)? \xnz.mem_r [453] : 
                        (N136)? \xnz.mem_r [486] : 
                        (N138)? \xnz.mem_r [519] : 
                        (N109)? \xnz.mem_r [552] : 
                        (N111)? \xnz.mem_r [585] : 
                        (N113)? \xnz.mem_r [618] : 
                        (N115)? \xnz.mem_r [651] : 
                        (N117)? \xnz.mem_r [684] : 
                        (N119)? \xnz.mem_r [717] : 
                        (N121)? \xnz.mem_r [750] : 
                        (N123)? \xnz.mem_r [783] : 
                        (N125)? \xnz.mem_r [816] : 
                        (N127)? \xnz.mem_r [849] : 
                        (N129)? \xnz.mem_r [882] : 
                        (N131)? \xnz.mem_r [915] : 
                        (N133)? \xnz.mem_r [948] : 
                        (N135)? \xnz.mem_r [981] : 
                        (N137)? \xnz.mem_r [1014] : 
                        (N139)? \xnz.mem_r [1047] : 1'b0;
  assign r_data_o[56] = (N108)? \xnz.mem_r [23] : 
                        (N110)? \xnz.mem_r [56] : 
                        (N112)? \xnz.mem_r [89] : 
                        (N114)? \xnz.mem_r [122] : 
                        (N116)? \xnz.mem_r [155] : 
                        (N118)? \xnz.mem_r [188] : 
                        (N120)? \xnz.mem_r [221] : 
                        (N122)? \xnz.mem_r [254] : 
                        (N124)? \xnz.mem_r [287] : 
                        (N126)? \xnz.mem_r [320] : 
                        (N128)? \xnz.mem_r [353] : 
                        (N130)? \xnz.mem_r [386] : 
                        (N132)? \xnz.mem_r [419] : 
                        (N134)? \xnz.mem_r [452] : 
                        (N136)? \xnz.mem_r [485] : 
                        (N138)? \xnz.mem_r [518] : 
                        (N109)? \xnz.mem_r [551] : 
                        (N111)? \xnz.mem_r [584] : 
                        (N113)? \xnz.mem_r [617] : 
                        (N115)? \xnz.mem_r [650] : 
                        (N117)? \xnz.mem_r [683] : 
                        (N119)? \xnz.mem_r [716] : 
                        (N121)? \xnz.mem_r [749] : 
                        (N123)? \xnz.mem_r [782] : 
                        (N125)? \xnz.mem_r [815] : 
                        (N127)? \xnz.mem_r [848] : 
                        (N129)? \xnz.mem_r [881] : 
                        (N131)? \xnz.mem_r [914] : 
                        (N133)? \xnz.mem_r [947] : 
                        (N135)? \xnz.mem_r [980] : 
                        (N137)? \xnz.mem_r [1013] : 
                        (N139)? \xnz.mem_r [1046] : 1'b0;
  assign r_data_o[55] = (N108)? \xnz.mem_r [22] : 
                        (N110)? \xnz.mem_r [55] : 
                        (N112)? \xnz.mem_r [88] : 
                        (N114)? \xnz.mem_r [121] : 
                        (N116)? \xnz.mem_r [154] : 
                        (N118)? \xnz.mem_r [187] : 
                        (N120)? \xnz.mem_r [220] : 
                        (N122)? \xnz.mem_r [253] : 
                        (N124)? \xnz.mem_r [286] : 
                        (N126)? \xnz.mem_r [319] : 
                        (N128)? \xnz.mem_r [352] : 
                        (N130)? \xnz.mem_r [385] : 
                        (N132)? \xnz.mem_r [418] : 
                        (N134)? \xnz.mem_r [451] : 
                        (N136)? \xnz.mem_r [484] : 
                        (N138)? \xnz.mem_r [517] : 
                        (N109)? \xnz.mem_r [550] : 
                        (N111)? \xnz.mem_r [583] : 
                        (N113)? \xnz.mem_r [616] : 
                        (N115)? \xnz.mem_r [649] : 
                        (N117)? \xnz.mem_r [682] : 
                        (N119)? \xnz.mem_r [715] : 
                        (N121)? \xnz.mem_r [748] : 
                        (N123)? \xnz.mem_r [781] : 
                        (N125)? \xnz.mem_r [814] : 
                        (N127)? \xnz.mem_r [847] : 
                        (N129)? \xnz.mem_r [880] : 
                        (N131)? \xnz.mem_r [913] : 
                        (N133)? \xnz.mem_r [946] : 
                        (N135)? \xnz.mem_r [979] : 
                        (N137)? \xnz.mem_r [1012] : 
                        (N139)? \xnz.mem_r [1045] : 1'b0;
  assign r_data_o[54] = (N108)? \xnz.mem_r [21] : 
                        (N110)? \xnz.mem_r [54] : 
                        (N112)? \xnz.mem_r [87] : 
                        (N114)? \xnz.mem_r [120] : 
                        (N116)? \xnz.mem_r [153] : 
                        (N118)? \xnz.mem_r [186] : 
                        (N120)? \xnz.mem_r [219] : 
                        (N122)? \xnz.mem_r [252] : 
                        (N124)? \xnz.mem_r [285] : 
                        (N126)? \xnz.mem_r [318] : 
                        (N128)? \xnz.mem_r [351] : 
                        (N130)? \xnz.mem_r [384] : 
                        (N132)? \xnz.mem_r [417] : 
                        (N134)? \xnz.mem_r [450] : 
                        (N136)? \xnz.mem_r [483] : 
                        (N138)? \xnz.mem_r [516] : 
                        (N109)? \xnz.mem_r [549] : 
                        (N111)? \xnz.mem_r [582] : 
                        (N113)? \xnz.mem_r [615] : 
                        (N115)? \xnz.mem_r [648] : 
                        (N117)? \xnz.mem_r [681] : 
                        (N119)? \xnz.mem_r [714] : 
                        (N121)? \xnz.mem_r [747] : 
                        (N123)? \xnz.mem_r [780] : 
                        (N125)? \xnz.mem_r [813] : 
                        (N127)? \xnz.mem_r [846] : 
                        (N129)? \xnz.mem_r [879] : 
                        (N131)? \xnz.mem_r [912] : 
                        (N133)? \xnz.mem_r [945] : 
                        (N135)? \xnz.mem_r [978] : 
                        (N137)? \xnz.mem_r [1011] : 
                        (N139)? \xnz.mem_r [1044] : 1'b0;
  assign r_data_o[53] = (N108)? \xnz.mem_r [20] : 
                        (N110)? \xnz.mem_r [53] : 
                        (N112)? \xnz.mem_r [86] : 
                        (N114)? \xnz.mem_r [119] : 
                        (N116)? \xnz.mem_r [152] : 
                        (N118)? \xnz.mem_r [185] : 
                        (N120)? \xnz.mem_r [218] : 
                        (N122)? \xnz.mem_r [251] : 
                        (N124)? \xnz.mem_r [284] : 
                        (N126)? \xnz.mem_r [317] : 
                        (N128)? \xnz.mem_r [350] : 
                        (N130)? \xnz.mem_r [383] : 
                        (N132)? \xnz.mem_r [416] : 
                        (N134)? \xnz.mem_r [449] : 
                        (N136)? \xnz.mem_r [482] : 
                        (N138)? \xnz.mem_r [515] : 
                        (N109)? \xnz.mem_r [548] : 
                        (N111)? \xnz.mem_r [581] : 
                        (N113)? \xnz.mem_r [614] : 
                        (N115)? \xnz.mem_r [647] : 
                        (N117)? \xnz.mem_r [680] : 
                        (N119)? \xnz.mem_r [713] : 
                        (N121)? \xnz.mem_r [746] : 
                        (N123)? \xnz.mem_r [779] : 
                        (N125)? \xnz.mem_r [812] : 
                        (N127)? \xnz.mem_r [845] : 
                        (N129)? \xnz.mem_r [878] : 
                        (N131)? \xnz.mem_r [911] : 
                        (N133)? \xnz.mem_r [944] : 
                        (N135)? \xnz.mem_r [977] : 
                        (N137)? \xnz.mem_r [1010] : 
                        (N139)? \xnz.mem_r [1043] : 1'b0;
  assign r_data_o[52] = (N108)? \xnz.mem_r [19] : 
                        (N110)? \xnz.mem_r [52] : 
                        (N112)? \xnz.mem_r [85] : 
                        (N114)? \xnz.mem_r [118] : 
                        (N116)? \xnz.mem_r [151] : 
                        (N118)? \xnz.mem_r [184] : 
                        (N120)? \xnz.mem_r [217] : 
                        (N122)? \xnz.mem_r [250] : 
                        (N124)? \xnz.mem_r [283] : 
                        (N126)? \xnz.mem_r [316] : 
                        (N128)? \xnz.mem_r [349] : 
                        (N130)? \xnz.mem_r [382] : 
                        (N132)? \xnz.mem_r [415] : 
                        (N134)? \xnz.mem_r [448] : 
                        (N136)? \xnz.mem_r [481] : 
                        (N138)? \xnz.mem_r [514] : 
                        (N109)? \xnz.mem_r [547] : 
                        (N111)? \xnz.mem_r [580] : 
                        (N113)? \xnz.mem_r [613] : 
                        (N115)? \xnz.mem_r [646] : 
                        (N117)? \xnz.mem_r [679] : 
                        (N119)? \xnz.mem_r [712] : 
                        (N121)? \xnz.mem_r [745] : 
                        (N123)? \xnz.mem_r [778] : 
                        (N125)? \xnz.mem_r [811] : 
                        (N127)? \xnz.mem_r [844] : 
                        (N129)? \xnz.mem_r [877] : 
                        (N131)? \xnz.mem_r [910] : 
                        (N133)? \xnz.mem_r [943] : 
                        (N135)? \xnz.mem_r [976] : 
                        (N137)? \xnz.mem_r [1009] : 
                        (N139)? \xnz.mem_r [1042] : 1'b0;
  assign r_data_o[51] = (N108)? \xnz.mem_r [18] : 
                        (N110)? \xnz.mem_r [51] : 
                        (N112)? \xnz.mem_r [84] : 
                        (N114)? \xnz.mem_r [117] : 
                        (N116)? \xnz.mem_r [150] : 
                        (N118)? \xnz.mem_r [183] : 
                        (N120)? \xnz.mem_r [216] : 
                        (N122)? \xnz.mem_r [249] : 
                        (N124)? \xnz.mem_r [282] : 
                        (N126)? \xnz.mem_r [315] : 
                        (N128)? \xnz.mem_r [348] : 
                        (N130)? \xnz.mem_r [381] : 
                        (N132)? \xnz.mem_r [414] : 
                        (N134)? \xnz.mem_r [447] : 
                        (N136)? \xnz.mem_r [480] : 
                        (N138)? \xnz.mem_r [513] : 
                        (N109)? \xnz.mem_r [546] : 
                        (N111)? \xnz.mem_r [579] : 
                        (N113)? \xnz.mem_r [612] : 
                        (N115)? \xnz.mem_r [645] : 
                        (N117)? \xnz.mem_r [678] : 
                        (N119)? \xnz.mem_r [711] : 
                        (N121)? \xnz.mem_r [744] : 
                        (N123)? \xnz.mem_r [777] : 
                        (N125)? \xnz.mem_r [810] : 
                        (N127)? \xnz.mem_r [843] : 
                        (N129)? \xnz.mem_r [876] : 
                        (N131)? \xnz.mem_r [909] : 
                        (N133)? \xnz.mem_r [942] : 
                        (N135)? \xnz.mem_r [975] : 
                        (N137)? \xnz.mem_r [1008] : 
                        (N139)? \xnz.mem_r [1041] : 1'b0;
  assign r_data_o[50] = (N108)? \xnz.mem_r [17] : 
                        (N110)? \xnz.mem_r [50] : 
                        (N112)? \xnz.mem_r [83] : 
                        (N114)? \xnz.mem_r [116] : 
                        (N116)? \xnz.mem_r [149] : 
                        (N118)? \xnz.mem_r [182] : 
                        (N120)? \xnz.mem_r [215] : 
                        (N122)? \xnz.mem_r [248] : 
                        (N124)? \xnz.mem_r [281] : 
                        (N126)? \xnz.mem_r [314] : 
                        (N128)? \xnz.mem_r [347] : 
                        (N130)? \xnz.mem_r [380] : 
                        (N132)? \xnz.mem_r [413] : 
                        (N134)? \xnz.mem_r [446] : 
                        (N136)? \xnz.mem_r [479] : 
                        (N138)? \xnz.mem_r [512] : 
                        (N109)? \xnz.mem_r [545] : 
                        (N111)? \xnz.mem_r [578] : 
                        (N113)? \xnz.mem_r [611] : 
                        (N115)? \xnz.mem_r [644] : 
                        (N117)? \xnz.mem_r [677] : 
                        (N119)? \xnz.mem_r [710] : 
                        (N121)? \xnz.mem_r [743] : 
                        (N123)? \xnz.mem_r [776] : 
                        (N125)? \xnz.mem_r [809] : 
                        (N127)? \xnz.mem_r [842] : 
                        (N129)? \xnz.mem_r [875] : 
                        (N131)? \xnz.mem_r [908] : 
                        (N133)? \xnz.mem_r [941] : 
                        (N135)? \xnz.mem_r [974] : 
                        (N137)? \xnz.mem_r [1007] : 
                        (N139)? \xnz.mem_r [1040] : 1'b0;
  assign r_data_o[49] = (N108)? \xnz.mem_r [16] : 
                        (N110)? \xnz.mem_r [49] : 
                        (N112)? \xnz.mem_r [82] : 
                        (N114)? \xnz.mem_r [115] : 
                        (N116)? \xnz.mem_r [148] : 
                        (N118)? \xnz.mem_r [181] : 
                        (N120)? \xnz.mem_r [214] : 
                        (N122)? \xnz.mem_r [247] : 
                        (N124)? \xnz.mem_r [280] : 
                        (N126)? \xnz.mem_r [313] : 
                        (N128)? \xnz.mem_r [346] : 
                        (N130)? \xnz.mem_r [379] : 
                        (N132)? \xnz.mem_r [412] : 
                        (N134)? \xnz.mem_r [445] : 
                        (N136)? \xnz.mem_r [478] : 
                        (N138)? \xnz.mem_r [511] : 
                        (N109)? \xnz.mem_r [544] : 
                        (N111)? \xnz.mem_r [577] : 
                        (N113)? \xnz.mem_r [610] : 
                        (N115)? \xnz.mem_r [643] : 
                        (N117)? \xnz.mem_r [676] : 
                        (N119)? \xnz.mem_r [709] : 
                        (N121)? \xnz.mem_r [742] : 
                        (N123)? \xnz.mem_r [775] : 
                        (N125)? \xnz.mem_r [808] : 
                        (N127)? \xnz.mem_r [841] : 
                        (N129)? \xnz.mem_r [874] : 
                        (N131)? \xnz.mem_r [907] : 
                        (N133)? \xnz.mem_r [940] : 
                        (N135)? \xnz.mem_r [973] : 
                        (N137)? \xnz.mem_r [1006] : 
                        (N139)? \xnz.mem_r [1039] : 1'b0;
  assign r_data_o[48] = (N108)? \xnz.mem_r [15] : 
                        (N110)? \xnz.mem_r [48] : 
                        (N112)? \xnz.mem_r [81] : 
                        (N114)? \xnz.mem_r [114] : 
                        (N116)? \xnz.mem_r [147] : 
                        (N118)? \xnz.mem_r [180] : 
                        (N120)? \xnz.mem_r [213] : 
                        (N122)? \xnz.mem_r [246] : 
                        (N124)? \xnz.mem_r [279] : 
                        (N126)? \xnz.mem_r [312] : 
                        (N128)? \xnz.mem_r [345] : 
                        (N130)? \xnz.mem_r [378] : 
                        (N132)? \xnz.mem_r [411] : 
                        (N134)? \xnz.mem_r [444] : 
                        (N136)? \xnz.mem_r [477] : 
                        (N138)? \xnz.mem_r [510] : 
                        (N109)? \xnz.mem_r [543] : 
                        (N111)? \xnz.mem_r [576] : 
                        (N113)? \xnz.mem_r [609] : 
                        (N115)? \xnz.mem_r [642] : 
                        (N117)? \xnz.mem_r [675] : 
                        (N119)? \xnz.mem_r [708] : 
                        (N121)? \xnz.mem_r [741] : 
                        (N123)? \xnz.mem_r [774] : 
                        (N125)? \xnz.mem_r [807] : 
                        (N127)? \xnz.mem_r [840] : 
                        (N129)? \xnz.mem_r [873] : 
                        (N131)? \xnz.mem_r [906] : 
                        (N133)? \xnz.mem_r [939] : 
                        (N135)? \xnz.mem_r [972] : 
                        (N137)? \xnz.mem_r [1005] : 
                        (N139)? \xnz.mem_r [1038] : 1'b0;
  assign r_data_o[47] = (N108)? \xnz.mem_r [14] : 
                        (N110)? \xnz.mem_r [47] : 
                        (N112)? \xnz.mem_r [80] : 
                        (N114)? \xnz.mem_r [113] : 
                        (N116)? \xnz.mem_r [146] : 
                        (N118)? \xnz.mem_r [179] : 
                        (N120)? \xnz.mem_r [212] : 
                        (N122)? \xnz.mem_r [245] : 
                        (N124)? \xnz.mem_r [278] : 
                        (N126)? \xnz.mem_r [311] : 
                        (N128)? \xnz.mem_r [344] : 
                        (N130)? \xnz.mem_r [377] : 
                        (N132)? \xnz.mem_r [410] : 
                        (N134)? \xnz.mem_r [443] : 
                        (N136)? \xnz.mem_r [476] : 
                        (N138)? \xnz.mem_r [509] : 
                        (N109)? \xnz.mem_r [542] : 
                        (N111)? \xnz.mem_r [575] : 
                        (N113)? \xnz.mem_r [608] : 
                        (N115)? \xnz.mem_r [641] : 
                        (N117)? \xnz.mem_r [674] : 
                        (N119)? \xnz.mem_r [707] : 
                        (N121)? \xnz.mem_r [740] : 
                        (N123)? \xnz.mem_r [773] : 
                        (N125)? \xnz.mem_r [806] : 
                        (N127)? \xnz.mem_r [839] : 
                        (N129)? \xnz.mem_r [872] : 
                        (N131)? \xnz.mem_r [905] : 
                        (N133)? \xnz.mem_r [938] : 
                        (N135)? \xnz.mem_r [971] : 
                        (N137)? \xnz.mem_r [1004] : 
                        (N139)? \xnz.mem_r [1037] : 1'b0;
  assign r_data_o[46] = (N108)? \xnz.mem_r [13] : 
                        (N110)? \xnz.mem_r [46] : 
                        (N112)? \xnz.mem_r [79] : 
                        (N114)? \xnz.mem_r [112] : 
                        (N116)? \xnz.mem_r [145] : 
                        (N118)? \xnz.mem_r [178] : 
                        (N120)? \xnz.mem_r [211] : 
                        (N122)? \xnz.mem_r [244] : 
                        (N124)? \xnz.mem_r [277] : 
                        (N126)? \xnz.mem_r [310] : 
                        (N128)? \xnz.mem_r [343] : 
                        (N130)? \xnz.mem_r [376] : 
                        (N132)? \xnz.mem_r [409] : 
                        (N134)? \xnz.mem_r [442] : 
                        (N136)? \xnz.mem_r [475] : 
                        (N138)? \xnz.mem_r [508] : 
                        (N109)? \xnz.mem_r [541] : 
                        (N111)? \xnz.mem_r [574] : 
                        (N113)? \xnz.mem_r [607] : 
                        (N115)? \xnz.mem_r [640] : 
                        (N117)? \xnz.mem_r [673] : 
                        (N119)? \xnz.mem_r [706] : 
                        (N121)? \xnz.mem_r [739] : 
                        (N123)? \xnz.mem_r [772] : 
                        (N125)? \xnz.mem_r [805] : 
                        (N127)? \xnz.mem_r [838] : 
                        (N129)? \xnz.mem_r [871] : 
                        (N131)? \xnz.mem_r [904] : 
                        (N133)? \xnz.mem_r [937] : 
                        (N135)? \xnz.mem_r [970] : 
                        (N137)? \xnz.mem_r [1003] : 
                        (N139)? \xnz.mem_r [1036] : 1'b0;
  assign r_data_o[45] = (N108)? \xnz.mem_r [12] : 
                        (N110)? \xnz.mem_r [45] : 
                        (N112)? \xnz.mem_r [78] : 
                        (N114)? \xnz.mem_r [111] : 
                        (N116)? \xnz.mem_r [144] : 
                        (N118)? \xnz.mem_r [177] : 
                        (N120)? \xnz.mem_r [210] : 
                        (N122)? \xnz.mem_r [243] : 
                        (N124)? \xnz.mem_r [276] : 
                        (N126)? \xnz.mem_r [309] : 
                        (N128)? \xnz.mem_r [342] : 
                        (N130)? \xnz.mem_r [375] : 
                        (N132)? \xnz.mem_r [408] : 
                        (N134)? \xnz.mem_r [441] : 
                        (N136)? \xnz.mem_r [474] : 
                        (N138)? \xnz.mem_r [507] : 
                        (N109)? \xnz.mem_r [540] : 
                        (N111)? \xnz.mem_r [573] : 
                        (N113)? \xnz.mem_r [606] : 
                        (N115)? \xnz.mem_r [639] : 
                        (N117)? \xnz.mem_r [672] : 
                        (N119)? \xnz.mem_r [705] : 
                        (N121)? \xnz.mem_r [738] : 
                        (N123)? \xnz.mem_r [771] : 
                        (N125)? \xnz.mem_r [804] : 
                        (N127)? \xnz.mem_r [837] : 
                        (N129)? \xnz.mem_r [870] : 
                        (N131)? \xnz.mem_r [903] : 
                        (N133)? \xnz.mem_r [936] : 
                        (N135)? \xnz.mem_r [969] : 
                        (N137)? \xnz.mem_r [1002] : 
                        (N139)? \xnz.mem_r [1035] : 1'b0;
  assign r_data_o[44] = (N108)? \xnz.mem_r [11] : 
                        (N110)? \xnz.mem_r [44] : 
                        (N112)? \xnz.mem_r [77] : 
                        (N114)? \xnz.mem_r [110] : 
                        (N116)? \xnz.mem_r [143] : 
                        (N118)? \xnz.mem_r [176] : 
                        (N120)? \xnz.mem_r [209] : 
                        (N122)? \xnz.mem_r [242] : 
                        (N124)? \xnz.mem_r [275] : 
                        (N126)? \xnz.mem_r [308] : 
                        (N128)? \xnz.mem_r [341] : 
                        (N130)? \xnz.mem_r [374] : 
                        (N132)? \xnz.mem_r [407] : 
                        (N134)? \xnz.mem_r [440] : 
                        (N136)? \xnz.mem_r [473] : 
                        (N138)? \xnz.mem_r [506] : 
                        (N109)? \xnz.mem_r [539] : 
                        (N111)? \xnz.mem_r [572] : 
                        (N113)? \xnz.mem_r [605] : 
                        (N115)? \xnz.mem_r [638] : 
                        (N117)? \xnz.mem_r [671] : 
                        (N119)? \xnz.mem_r [704] : 
                        (N121)? \xnz.mem_r [737] : 
                        (N123)? \xnz.mem_r [770] : 
                        (N125)? \xnz.mem_r [803] : 
                        (N127)? \xnz.mem_r [836] : 
                        (N129)? \xnz.mem_r [869] : 
                        (N131)? \xnz.mem_r [902] : 
                        (N133)? \xnz.mem_r [935] : 
                        (N135)? \xnz.mem_r [968] : 
                        (N137)? \xnz.mem_r [1001] : 
                        (N139)? \xnz.mem_r [1034] : 1'b0;
  assign r_data_o[43] = (N108)? \xnz.mem_r [10] : 
                        (N110)? \xnz.mem_r [43] : 
                        (N112)? \xnz.mem_r [76] : 
                        (N114)? \xnz.mem_r [109] : 
                        (N116)? \xnz.mem_r [142] : 
                        (N118)? \xnz.mem_r [175] : 
                        (N120)? \xnz.mem_r [208] : 
                        (N122)? \xnz.mem_r [241] : 
                        (N124)? \xnz.mem_r [274] : 
                        (N126)? \xnz.mem_r [307] : 
                        (N128)? \xnz.mem_r [340] : 
                        (N130)? \xnz.mem_r [373] : 
                        (N132)? \xnz.mem_r [406] : 
                        (N134)? \xnz.mem_r [439] : 
                        (N136)? \xnz.mem_r [472] : 
                        (N138)? \xnz.mem_r [505] : 
                        (N109)? \xnz.mem_r [538] : 
                        (N111)? \xnz.mem_r [571] : 
                        (N113)? \xnz.mem_r [604] : 
                        (N115)? \xnz.mem_r [637] : 
                        (N117)? \xnz.mem_r [670] : 
                        (N119)? \xnz.mem_r [703] : 
                        (N121)? \xnz.mem_r [736] : 
                        (N123)? \xnz.mem_r [769] : 
                        (N125)? \xnz.mem_r [802] : 
                        (N127)? \xnz.mem_r [835] : 
                        (N129)? \xnz.mem_r [868] : 
                        (N131)? \xnz.mem_r [901] : 
                        (N133)? \xnz.mem_r [934] : 
                        (N135)? \xnz.mem_r [967] : 
                        (N137)? \xnz.mem_r [1000] : 
                        (N139)? \xnz.mem_r [1033] : 1'b0;
  assign r_data_o[42] = (N108)? \xnz.mem_r [9] : 
                        (N110)? \xnz.mem_r [42] : 
                        (N112)? \xnz.mem_r [75] : 
                        (N114)? \xnz.mem_r [108] : 
                        (N116)? \xnz.mem_r [141] : 
                        (N118)? \xnz.mem_r [174] : 
                        (N120)? \xnz.mem_r [207] : 
                        (N122)? \xnz.mem_r [240] : 
                        (N124)? \xnz.mem_r [273] : 
                        (N126)? \xnz.mem_r [306] : 
                        (N128)? \xnz.mem_r [339] : 
                        (N130)? \xnz.mem_r [372] : 
                        (N132)? \xnz.mem_r [405] : 
                        (N134)? \xnz.mem_r [438] : 
                        (N136)? \xnz.mem_r [471] : 
                        (N138)? \xnz.mem_r [504] : 
                        (N109)? \xnz.mem_r [537] : 
                        (N111)? \xnz.mem_r [570] : 
                        (N113)? \xnz.mem_r [603] : 
                        (N115)? \xnz.mem_r [636] : 
                        (N117)? \xnz.mem_r [669] : 
                        (N119)? \xnz.mem_r [702] : 
                        (N121)? \xnz.mem_r [735] : 
                        (N123)? \xnz.mem_r [768] : 
                        (N125)? \xnz.mem_r [801] : 
                        (N127)? \xnz.mem_r [834] : 
                        (N129)? \xnz.mem_r [867] : 
                        (N131)? \xnz.mem_r [900] : 
                        (N133)? \xnz.mem_r [933] : 
                        (N135)? \xnz.mem_r [966] : 
                        (N137)? \xnz.mem_r [999] : 
                        (N139)? \xnz.mem_r [1032] : 1'b0;
  assign r_data_o[41] = (N108)? \xnz.mem_r [8] : 
                        (N110)? \xnz.mem_r [41] : 
                        (N112)? \xnz.mem_r [74] : 
                        (N114)? \xnz.mem_r [107] : 
                        (N116)? \xnz.mem_r [140] : 
                        (N118)? \xnz.mem_r [173] : 
                        (N120)? \xnz.mem_r [206] : 
                        (N122)? \xnz.mem_r [239] : 
                        (N124)? \xnz.mem_r [272] : 
                        (N126)? \xnz.mem_r [305] : 
                        (N128)? \xnz.mem_r [338] : 
                        (N130)? \xnz.mem_r [371] : 
                        (N132)? \xnz.mem_r [404] : 
                        (N134)? \xnz.mem_r [437] : 
                        (N136)? \xnz.mem_r [470] : 
                        (N138)? \xnz.mem_r [503] : 
                        (N109)? \xnz.mem_r [536] : 
                        (N111)? \xnz.mem_r [569] : 
                        (N113)? \xnz.mem_r [602] : 
                        (N115)? \xnz.mem_r [635] : 
                        (N117)? \xnz.mem_r [668] : 
                        (N119)? \xnz.mem_r [701] : 
                        (N121)? \xnz.mem_r [734] : 
                        (N123)? \xnz.mem_r [767] : 
                        (N125)? \xnz.mem_r [800] : 
                        (N127)? \xnz.mem_r [833] : 
                        (N129)? \xnz.mem_r [866] : 
                        (N131)? \xnz.mem_r [899] : 
                        (N133)? \xnz.mem_r [932] : 
                        (N135)? \xnz.mem_r [965] : 
                        (N137)? \xnz.mem_r [998] : 
                        (N139)? \xnz.mem_r [1031] : 1'b0;
  assign r_data_o[40] = (N108)? \xnz.mem_r [7] : 
                        (N110)? \xnz.mem_r [40] : 
                        (N112)? \xnz.mem_r [73] : 
                        (N114)? \xnz.mem_r [106] : 
                        (N116)? \xnz.mem_r [139] : 
                        (N118)? \xnz.mem_r [172] : 
                        (N120)? \xnz.mem_r [205] : 
                        (N122)? \xnz.mem_r [238] : 
                        (N124)? \xnz.mem_r [271] : 
                        (N126)? \xnz.mem_r [304] : 
                        (N128)? \xnz.mem_r [337] : 
                        (N130)? \xnz.mem_r [370] : 
                        (N132)? \xnz.mem_r [403] : 
                        (N134)? \xnz.mem_r [436] : 
                        (N136)? \xnz.mem_r [469] : 
                        (N138)? \xnz.mem_r [502] : 
                        (N109)? \xnz.mem_r [535] : 
                        (N111)? \xnz.mem_r [568] : 
                        (N113)? \xnz.mem_r [601] : 
                        (N115)? \xnz.mem_r [634] : 
                        (N117)? \xnz.mem_r [667] : 
                        (N119)? \xnz.mem_r [700] : 
                        (N121)? \xnz.mem_r [733] : 
                        (N123)? \xnz.mem_r [766] : 
                        (N125)? \xnz.mem_r [799] : 
                        (N127)? \xnz.mem_r [832] : 
                        (N129)? \xnz.mem_r [865] : 
                        (N131)? \xnz.mem_r [898] : 
                        (N133)? \xnz.mem_r [931] : 
                        (N135)? \xnz.mem_r [964] : 
                        (N137)? \xnz.mem_r [997] : 
                        (N139)? \xnz.mem_r [1030] : 1'b0;
  assign r_data_o[39] = (N108)? \xnz.mem_r [6] : 
                        (N110)? \xnz.mem_r [39] : 
                        (N112)? \xnz.mem_r [72] : 
                        (N114)? \xnz.mem_r [105] : 
                        (N116)? \xnz.mem_r [138] : 
                        (N118)? \xnz.mem_r [171] : 
                        (N120)? \xnz.mem_r [204] : 
                        (N122)? \xnz.mem_r [237] : 
                        (N124)? \xnz.mem_r [270] : 
                        (N126)? \xnz.mem_r [303] : 
                        (N128)? \xnz.mem_r [336] : 
                        (N130)? \xnz.mem_r [369] : 
                        (N132)? \xnz.mem_r [402] : 
                        (N134)? \xnz.mem_r [435] : 
                        (N136)? \xnz.mem_r [468] : 
                        (N138)? \xnz.mem_r [501] : 
                        (N109)? \xnz.mem_r [534] : 
                        (N111)? \xnz.mem_r [567] : 
                        (N113)? \xnz.mem_r [600] : 
                        (N115)? \xnz.mem_r [633] : 
                        (N117)? \xnz.mem_r [666] : 
                        (N119)? \xnz.mem_r [699] : 
                        (N121)? \xnz.mem_r [732] : 
                        (N123)? \xnz.mem_r [765] : 
                        (N125)? \xnz.mem_r [798] : 
                        (N127)? \xnz.mem_r [831] : 
                        (N129)? \xnz.mem_r [864] : 
                        (N131)? \xnz.mem_r [897] : 
                        (N133)? \xnz.mem_r [930] : 
                        (N135)? \xnz.mem_r [963] : 
                        (N137)? \xnz.mem_r [996] : 
                        (N139)? \xnz.mem_r [1029] : 1'b0;
  assign r_data_o[38] = (N108)? \xnz.mem_r [5] : 
                        (N110)? \xnz.mem_r [38] : 
                        (N112)? \xnz.mem_r [71] : 
                        (N114)? \xnz.mem_r [104] : 
                        (N116)? \xnz.mem_r [137] : 
                        (N118)? \xnz.mem_r [170] : 
                        (N120)? \xnz.mem_r [203] : 
                        (N122)? \xnz.mem_r [236] : 
                        (N124)? \xnz.mem_r [269] : 
                        (N126)? \xnz.mem_r [302] : 
                        (N128)? \xnz.mem_r [335] : 
                        (N130)? \xnz.mem_r [368] : 
                        (N132)? \xnz.mem_r [401] : 
                        (N134)? \xnz.mem_r [434] : 
                        (N136)? \xnz.mem_r [467] : 
                        (N138)? \xnz.mem_r [500] : 
                        (N109)? \xnz.mem_r [533] : 
                        (N111)? \xnz.mem_r [566] : 
                        (N113)? \xnz.mem_r [599] : 
                        (N115)? \xnz.mem_r [632] : 
                        (N117)? \xnz.mem_r [665] : 
                        (N119)? \xnz.mem_r [698] : 
                        (N121)? \xnz.mem_r [731] : 
                        (N123)? \xnz.mem_r [764] : 
                        (N125)? \xnz.mem_r [797] : 
                        (N127)? \xnz.mem_r [830] : 
                        (N129)? \xnz.mem_r [863] : 
                        (N131)? \xnz.mem_r [896] : 
                        (N133)? \xnz.mem_r [929] : 
                        (N135)? \xnz.mem_r [962] : 
                        (N137)? \xnz.mem_r [995] : 
                        (N139)? \xnz.mem_r [1028] : 1'b0;
  assign r_data_o[37] = (N108)? \xnz.mem_r [4] : 
                        (N110)? \xnz.mem_r [37] : 
                        (N112)? \xnz.mem_r [70] : 
                        (N114)? \xnz.mem_r [103] : 
                        (N116)? \xnz.mem_r [136] : 
                        (N118)? \xnz.mem_r [169] : 
                        (N120)? \xnz.mem_r [202] : 
                        (N122)? \xnz.mem_r [235] : 
                        (N124)? \xnz.mem_r [268] : 
                        (N126)? \xnz.mem_r [301] : 
                        (N128)? \xnz.mem_r [334] : 
                        (N130)? \xnz.mem_r [367] : 
                        (N132)? \xnz.mem_r [400] : 
                        (N134)? \xnz.mem_r [433] : 
                        (N136)? \xnz.mem_r [466] : 
                        (N138)? \xnz.mem_r [499] : 
                        (N109)? \xnz.mem_r [532] : 
                        (N111)? \xnz.mem_r [565] : 
                        (N113)? \xnz.mem_r [598] : 
                        (N115)? \xnz.mem_r [631] : 
                        (N117)? \xnz.mem_r [664] : 
                        (N119)? \xnz.mem_r [697] : 
                        (N121)? \xnz.mem_r [730] : 
                        (N123)? \xnz.mem_r [763] : 
                        (N125)? \xnz.mem_r [796] : 
                        (N127)? \xnz.mem_r [829] : 
                        (N129)? \xnz.mem_r [862] : 
                        (N131)? \xnz.mem_r [895] : 
                        (N133)? \xnz.mem_r [928] : 
                        (N135)? \xnz.mem_r [961] : 
                        (N137)? \xnz.mem_r [994] : 
                        (N139)? \xnz.mem_r [1027] : 1'b0;
  assign r_data_o[36] = (N108)? \xnz.mem_r [3] : 
                        (N110)? \xnz.mem_r [36] : 
                        (N112)? \xnz.mem_r [69] : 
                        (N114)? \xnz.mem_r [102] : 
                        (N116)? \xnz.mem_r [135] : 
                        (N118)? \xnz.mem_r [168] : 
                        (N120)? \xnz.mem_r [201] : 
                        (N122)? \xnz.mem_r [234] : 
                        (N124)? \xnz.mem_r [267] : 
                        (N126)? \xnz.mem_r [300] : 
                        (N128)? \xnz.mem_r [333] : 
                        (N130)? \xnz.mem_r [366] : 
                        (N132)? \xnz.mem_r [399] : 
                        (N134)? \xnz.mem_r [432] : 
                        (N136)? \xnz.mem_r [465] : 
                        (N138)? \xnz.mem_r [498] : 
                        (N109)? \xnz.mem_r [531] : 
                        (N111)? \xnz.mem_r [564] : 
                        (N113)? \xnz.mem_r [597] : 
                        (N115)? \xnz.mem_r [630] : 
                        (N117)? \xnz.mem_r [663] : 
                        (N119)? \xnz.mem_r [696] : 
                        (N121)? \xnz.mem_r [729] : 
                        (N123)? \xnz.mem_r [762] : 
                        (N125)? \xnz.mem_r [795] : 
                        (N127)? \xnz.mem_r [828] : 
                        (N129)? \xnz.mem_r [861] : 
                        (N131)? \xnz.mem_r [894] : 
                        (N133)? \xnz.mem_r [927] : 
                        (N135)? \xnz.mem_r [960] : 
                        (N137)? \xnz.mem_r [993] : 
                        (N139)? \xnz.mem_r [1026] : 1'b0;
  assign r_data_o[35] = (N108)? \xnz.mem_r [2] : 
                        (N110)? \xnz.mem_r [35] : 
                        (N112)? \xnz.mem_r [68] : 
                        (N114)? \xnz.mem_r [101] : 
                        (N116)? \xnz.mem_r [134] : 
                        (N118)? \xnz.mem_r [167] : 
                        (N120)? \xnz.mem_r [200] : 
                        (N122)? \xnz.mem_r [233] : 
                        (N124)? \xnz.mem_r [266] : 
                        (N126)? \xnz.mem_r [299] : 
                        (N128)? \xnz.mem_r [332] : 
                        (N130)? \xnz.mem_r [365] : 
                        (N132)? \xnz.mem_r [398] : 
                        (N134)? \xnz.mem_r [431] : 
                        (N136)? \xnz.mem_r [464] : 
                        (N138)? \xnz.mem_r [497] : 
                        (N109)? \xnz.mem_r [530] : 
                        (N111)? \xnz.mem_r [563] : 
                        (N113)? \xnz.mem_r [596] : 
                        (N115)? \xnz.mem_r [629] : 
                        (N117)? \xnz.mem_r [662] : 
                        (N119)? \xnz.mem_r [695] : 
                        (N121)? \xnz.mem_r [728] : 
                        (N123)? \xnz.mem_r [761] : 
                        (N125)? \xnz.mem_r [794] : 
                        (N127)? \xnz.mem_r [827] : 
                        (N129)? \xnz.mem_r [860] : 
                        (N131)? \xnz.mem_r [893] : 
                        (N133)? \xnz.mem_r [926] : 
                        (N135)? \xnz.mem_r [959] : 
                        (N137)? \xnz.mem_r [992] : 
                        (N139)? \xnz.mem_r [1025] : 1'b0;
  assign r_data_o[34] = (N108)? \xnz.mem_r [1] : 
                        (N110)? \xnz.mem_r [34] : 
                        (N112)? \xnz.mem_r [67] : 
                        (N114)? \xnz.mem_r [100] : 
                        (N116)? \xnz.mem_r [133] : 
                        (N118)? \xnz.mem_r [166] : 
                        (N120)? \xnz.mem_r [199] : 
                        (N122)? \xnz.mem_r [232] : 
                        (N124)? \xnz.mem_r [265] : 
                        (N126)? \xnz.mem_r [298] : 
                        (N128)? \xnz.mem_r [331] : 
                        (N130)? \xnz.mem_r [364] : 
                        (N132)? \xnz.mem_r [397] : 
                        (N134)? \xnz.mem_r [430] : 
                        (N136)? \xnz.mem_r [463] : 
                        (N138)? \xnz.mem_r [496] : 
                        (N109)? \xnz.mem_r [529] : 
                        (N111)? \xnz.mem_r [562] : 
                        (N113)? \xnz.mem_r [595] : 
                        (N115)? \xnz.mem_r [628] : 
                        (N117)? \xnz.mem_r [661] : 
                        (N119)? \xnz.mem_r [694] : 
                        (N121)? \xnz.mem_r [727] : 
                        (N123)? \xnz.mem_r [760] : 
                        (N125)? \xnz.mem_r [793] : 
                        (N127)? \xnz.mem_r [826] : 
                        (N129)? \xnz.mem_r [859] : 
                        (N131)? \xnz.mem_r [892] : 
                        (N133)? \xnz.mem_r [925] : 
                        (N135)? \xnz.mem_r [958] : 
                        (N137)? \xnz.mem_r [991] : 
                        (N139)? \xnz.mem_r [1024] : 1'b0;
  assign r_data_o[33] = (N108)? \xnz.mem_r [0] : 
                        (N110)? \xnz.mem_r [33] : 
                        (N112)? \xnz.mem_r [66] : 
                        (N114)? \xnz.mem_r [99] : 
                        (N116)? \xnz.mem_r [132] : 
                        (N118)? \xnz.mem_r [165] : 
                        (N120)? \xnz.mem_r [198] : 
                        (N122)? \xnz.mem_r [231] : 
                        (N124)? \xnz.mem_r [264] : 
                        (N126)? \xnz.mem_r [297] : 
                        (N128)? \xnz.mem_r [330] : 
                        (N130)? \xnz.mem_r [363] : 
                        (N132)? \xnz.mem_r [396] : 
                        (N134)? \xnz.mem_r [429] : 
                        (N136)? \xnz.mem_r [462] : 
                        (N138)? \xnz.mem_r [495] : 
                        (N109)? \xnz.mem_r [528] : 
                        (N111)? \xnz.mem_r [561] : 
                        (N113)? \xnz.mem_r [594] : 
                        (N115)? \xnz.mem_r [627] : 
                        (N117)? \xnz.mem_r [660] : 
                        (N119)? \xnz.mem_r [693] : 
                        (N121)? \xnz.mem_r [726] : 
                        (N123)? \xnz.mem_r [759] : 
                        (N125)? \xnz.mem_r [792] : 
                        (N127)? \xnz.mem_r [825] : 
                        (N129)? \xnz.mem_r [858] : 
                        (N131)? \xnz.mem_r [891] : 
                        (N133)? \xnz.mem_r [924] : 
                        (N135)? \xnz.mem_r [957] : 
                        (N137)? \xnz.mem_r [990] : 
                        (N139)? \xnz.mem_r [1023] : 1'b0;
  assign r_data_o[98] = (N173)? \xnz.mem_r [32] : 
                        (N175)? \xnz.mem_r [65] : 
                        (N177)? \xnz.mem_r [98] : 
                        (N179)? \xnz.mem_r [131] : 
                        (N181)? \xnz.mem_r [164] : 
                        (N183)? \xnz.mem_r [197] : 
                        (N185)? \xnz.mem_r [230] : 
                        (N187)? \xnz.mem_r [263] : 
                        (N189)? \xnz.mem_r [296] : 
                        (N191)? \xnz.mem_r [329] : 
                        (N193)? \xnz.mem_r [362] : 
                        (N195)? \xnz.mem_r [395] : 
                        (N197)? \xnz.mem_r [428] : 
                        (N199)? \xnz.mem_r [461] : 
                        (N201)? \xnz.mem_r [494] : 
                        (N203)? \xnz.mem_r [527] : 
                        (N174)? \xnz.mem_r [560] : 
                        (N176)? \xnz.mem_r [593] : 
                        (N178)? \xnz.mem_r [626] : 
                        (N180)? \xnz.mem_r [659] : 
                        (N182)? \xnz.mem_r [692] : 
                        (N184)? \xnz.mem_r [725] : 
                        (N186)? \xnz.mem_r [758] : 
                        (N188)? \xnz.mem_r [791] : 
                        (N190)? \xnz.mem_r [824] : 
                        (N192)? \xnz.mem_r [857] : 
                        (N194)? \xnz.mem_r [890] : 
                        (N196)? \xnz.mem_r [923] : 
                        (N198)? \xnz.mem_r [956] : 
                        (N200)? \xnz.mem_r [989] : 
                        (N202)? \xnz.mem_r [1022] : 
                        (N204)? \xnz.mem_r [1055] : 1'b0;
  assign r_data_o[97] = (N173)? \xnz.mem_r [31] : 
                        (N175)? \xnz.mem_r [64] : 
                        (N177)? \xnz.mem_r [97] : 
                        (N179)? \xnz.mem_r [130] : 
                        (N181)? \xnz.mem_r [163] : 
                        (N183)? \xnz.mem_r [196] : 
                        (N185)? \xnz.mem_r [229] : 
                        (N187)? \xnz.mem_r [262] : 
                        (N189)? \xnz.mem_r [295] : 
                        (N191)? \xnz.mem_r [328] : 
                        (N193)? \xnz.mem_r [361] : 
                        (N195)? \xnz.mem_r [394] : 
                        (N197)? \xnz.mem_r [427] : 
                        (N199)? \xnz.mem_r [460] : 
                        (N201)? \xnz.mem_r [493] : 
                        (N203)? \xnz.mem_r [526] : 
                        (N174)? \xnz.mem_r [559] : 
                        (N176)? \xnz.mem_r [592] : 
                        (N178)? \xnz.mem_r [625] : 
                        (N180)? \xnz.mem_r [658] : 
                        (N182)? \xnz.mem_r [691] : 
                        (N184)? \xnz.mem_r [724] : 
                        (N186)? \xnz.mem_r [757] : 
                        (N188)? \xnz.mem_r [790] : 
                        (N190)? \xnz.mem_r [823] : 
                        (N192)? \xnz.mem_r [856] : 
                        (N194)? \xnz.mem_r [889] : 
                        (N196)? \xnz.mem_r [922] : 
                        (N198)? \xnz.mem_r [955] : 
                        (N200)? \xnz.mem_r [988] : 
                        (N202)? \xnz.mem_r [1021] : 
                        (N204)? \xnz.mem_r [1054] : 1'b0;
  assign r_data_o[96] = (N173)? \xnz.mem_r [30] : 
                        (N175)? \xnz.mem_r [63] : 
                        (N177)? \xnz.mem_r [96] : 
                        (N179)? \xnz.mem_r [129] : 
                        (N181)? \xnz.mem_r [162] : 
                        (N183)? \xnz.mem_r [195] : 
                        (N185)? \xnz.mem_r [228] : 
                        (N187)? \xnz.mem_r [261] : 
                        (N189)? \xnz.mem_r [294] : 
                        (N191)? \xnz.mem_r [327] : 
                        (N193)? \xnz.mem_r [360] : 
                        (N195)? \xnz.mem_r [393] : 
                        (N197)? \xnz.mem_r [426] : 
                        (N199)? \xnz.mem_r [459] : 
                        (N201)? \xnz.mem_r [492] : 
                        (N203)? \xnz.mem_r [525] : 
                        (N174)? \xnz.mem_r [558] : 
                        (N176)? \xnz.mem_r [591] : 
                        (N178)? \xnz.mem_r [624] : 
                        (N180)? \xnz.mem_r [657] : 
                        (N182)? \xnz.mem_r [690] : 
                        (N184)? \xnz.mem_r [723] : 
                        (N186)? \xnz.mem_r [756] : 
                        (N188)? \xnz.mem_r [789] : 
                        (N190)? \xnz.mem_r [822] : 
                        (N192)? \xnz.mem_r [855] : 
                        (N194)? \xnz.mem_r [888] : 
                        (N196)? \xnz.mem_r [921] : 
                        (N198)? \xnz.mem_r [954] : 
                        (N200)? \xnz.mem_r [987] : 
                        (N202)? \xnz.mem_r [1020] : 
                        (N204)? \xnz.mem_r [1053] : 1'b0;
  assign r_data_o[95] = (N173)? \xnz.mem_r [29] : 
                        (N175)? \xnz.mem_r [62] : 
                        (N177)? \xnz.mem_r [95] : 
                        (N179)? \xnz.mem_r [128] : 
                        (N181)? \xnz.mem_r [161] : 
                        (N183)? \xnz.mem_r [194] : 
                        (N185)? \xnz.mem_r [227] : 
                        (N187)? \xnz.mem_r [260] : 
                        (N189)? \xnz.mem_r [293] : 
                        (N191)? \xnz.mem_r [326] : 
                        (N193)? \xnz.mem_r [359] : 
                        (N195)? \xnz.mem_r [392] : 
                        (N197)? \xnz.mem_r [425] : 
                        (N199)? \xnz.mem_r [458] : 
                        (N201)? \xnz.mem_r [491] : 
                        (N203)? \xnz.mem_r [524] : 
                        (N174)? \xnz.mem_r [557] : 
                        (N176)? \xnz.mem_r [590] : 
                        (N178)? \xnz.mem_r [623] : 
                        (N180)? \xnz.mem_r [656] : 
                        (N182)? \xnz.mem_r [689] : 
                        (N184)? \xnz.mem_r [722] : 
                        (N186)? \xnz.mem_r [755] : 
                        (N188)? \xnz.mem_r [788] : 
                        (N190)? \xnz.mem_r [821] : 
                        (N192)? \xnz.mem_r [854] : 
                        (N194)? \xnz.mem_r [887] : 
                        (N196)? \xnz.mem_r [920] : 
                        (N198)? \xnz.mem_r [953] : 
                        (N200)? \xnz.mem_r [986] : 
                        (N202)? \xnz.mem_r [1019] : 
                        (N204)? \xnz.mem_r [1052] : 1'b0;
  assign r_data_o[94] = (N173)? \xnz.mem_r [28] : 
                        (N175)? \xnz.mem_r [61] : 
                        (N177)? \xnz.mem_r [94] : 
                        (N179)? \xnz.mem_r [127] : 
                        (N181)? \xnz.mem_r [160] : 
                        (N183)? \xnz.mem_r [193] : 
                        (N185)? \xnz.mem_r [226] : 
                        (N187)? \xnz.mem_r [259] : 
                        (N189)? \xnz.mem_r [292] : 
                        (N191)? \xnz.mem_r [325] : 
                        (N193)? \xnz.mem_r [358] : 
                        (N195)? \xnz.mem_r [391] : 
                        (N197)? \xnz.mem_r [424] : 
                        (N199)? \xnz.mem_r [457] : 
                        (N201)? \xnz.mem_r [490] : 
                        (N203)? \xnz.mem_r [523] : 
                        (N174)? \xnz.mem_r [556] : 
                        (N176)? \xnz.mem_r [589] : 
                        (N178)? \xnz.mem_r [622] : 
                        (N180)? \xnz.mem_r [655] : 
                        (N182)? \xnz.mem_r [688] : 
                        (N184)? \xnz.mem_r [721] : 
                        (N186)? \xnz.mem_r [754] : 
                        (N188)? \xnz.mem_r [787] : 
                        (N190)? \xnz.mem_r [820] : 
                        (N192)? \xnz.mem_r [853] : 
                        (N194)? \xnz.mem_r [886] : 
                        (N196)? \xnz.mem_r [919] : 
                        (N198)? \xnz.mem_r [952] : 
                        (N200)? \xnz.mem_r [985] : 
                        (N202)? \xnz.mem_r [1018] : 
                        (N204)? \xnz.mem_r [1051] : 1'b0;
  assign r_data_o[93] = (N173)? \xnz.mem_r [27] : 
                        (N175)? \xnz.mem_r [60] : 
                        (N177)? \xnz.mem_r [93] : 
                        (N179)? \xnz.mem_r [126] : 
                        (N181)? \xnz.mem_r [159] : 
                        (N183)? \xnz.mem_r [192] : 
                        (N185)? \xnz.mem_r [225] : 
                        (N187)? \xnz.mem_r [258] : 
                        (N189)? \xnz.mem_r [291] : 
                        (N191)? \xnz.mem_r [324] : 
                        (N193)? \xnz.mem_r [357] : 
                        (N195)? \xnz.mem_r [390] : 
                        (N197)? \xnz.mem_r [423] : 
                        (N199)? \xnz.mem_r [456] : 
                        (N201)? \xnz.mem_r [489] : 
                        (N203)? \xnz.mem_r [522] : 
                        (N174)? \xnz.mem_r [555] : 
                        (N176)? \xnz.mem_r [588] : 
                        (N178)? \xnz.mem_r [621] : 
                        (N180)? \xnz.mem_r [654] : 
                        (N182)? \xnz.mem_r [687] : 
                        (N184)? \xnz.mem_r [720] : 
                        (N186)? \xnz.mem_r [753] : 
                        (N188)? \xnz.mem_r [786] : 
                        (N190)? \xnz.mem_r [819] : 
                        (N192)? \xnz.mem_r [852] : 
                        (N194)? \xnz.mem_r [885] : 
                        (N196)? \xnz.mem_r [918] : 
                        (N198)? \xnz.mem_r [951] : 
                        (N200)? \xnz.mem_r [984] : 
                        (N202)? \xnz.mem_r [1017] : 
                        (N204)? \xnz.mem_r [1050] : 1'b0;
  assign r_data_o[92] = (N173)? \xnz.mem_r [26] : 
                        (N175)? \xnz.mem_r [59] : 
                        (N177)? \xnz.mem_r [92] : 
                        (N179)? \xnz.mem_r [125] : 
                        (N181)? \xnz.mem_r [158] : 
                        (N183)? \xnz.mem_r [191] : 
                        (N185)? \xnz.mem_r [224] : 
                        (N187)? \xnz.mem_r [257] : 
                        (N189)? \xnz.mem_r [290] : 
                        (N191)? \xnz.mem_r [323] : 
                        (N193)? \xnz.mem_r [356] : 
                        (N195)? \xnz.mem_r [389] : 
                        (N197)? \xnz.mem_r [422] : 
                        (N199)? \xnz.mem_r [455] : 
                        (N201)? \xnz.mem_r [488] : 
                        (N203)? \xnz.mem_r [521] : 
                        (N174)? \xnz.mem_r [554] : 
                        (N176)? \xnz.mem_r [587] : 
                        (N178)? \xnz.mem_r [620] : 
                        (N180)? \xnz.mem_r [653] : 
                        (N182)? \xnz.mem_r [686] : 
                        (N184)? \xnz.mem_r [719] : 
                        (N186)? \xnz.mem_r [752] : 
                        (N188)? \xnz.mem_r [785] : 
                        (N190)? \xnz.mem_r [818] : 
                        (N192)? \xnz.mem_r [851] : 
                        (N194)? \xnz.mem_r [884] : 
                        (N196)? \xnz.mem_r [917] : 
                        (N198)? \xnz.mem_r [950] : 
                        (N200)? \xnz.mem_r [983] : 
                        (N202)? \xnz.mem_r [1016] : 
                        (N204)? \xnz.mem_r [1049] : 1'b0;
  assign r_data_o[91] = (N173)? \xnz.mem_r [25] : 
                        (N175)? \xnz.mem_r [58] : 
                        (N177)? \xnz.mem_r [91] : 
                        (N179)? \xnz.mem_r [124] : 
                        (N181)? \xnz.mem_r [157] : 
                        (N183)? \xnz.mem_r [190] : 
                        (N185)? \xnz.mem_r [223] : 
                        (N187)? \xnz.mem_r [256] : 
                        (N189)? \xnz.mem_r [289] : 
                        (N191)? \xnz.mem_r [322] : 
                        (N193)? \xnz.mem_r [355] : 
                        (N195)? \xnz.mem_r [388] : 
                        (N197)? \xnz.mem_r [421] : 
                        (N199)? \xnz.mem_r [454] : 
                        (N201)? \xnz.mem_r [487] : 
                        (N203)? \xnz.mem_r [520] : 
                        (N174)? \xnz.mem_r [553] : 
                        (N176)? \xnz.mem_r [586] : 
                        (N178)? \xnz.mem_r [619] : 
                        (N180)? \xnz.mem_r [652] : 
                        (N182)? \xnz.mem_r [685] : 
                        (N184)? \xnz.mem_r [718] : 
                        (N186)? \xnz.mem_r [751] : 
                        (N188)? \xnz.mem_r [784] : 
                        (N190)? \xnz.mem_r [817] : 
                        (N192)? \xnz.mem_r [850] : 
                        (N194)? \xnz.mem_r [883] : 
                        (N196)? \xnz.mem_r [916] : 
                        (N198)? \xnz.mem_r [949] : 
                        (N200)? \xnz.mem_r [982] : 
                        (N202)? \xnz.mem_r [1015] : 
                        (N204)? \xnz.mem_r [1048] : 1'b0;
  assign r_data_o[90] = (N173)? \xnz.mem_r [24] : 
                        (N175)? \xnz.mem_r [57] : 
                        (N177)? \xnz.mem_r [90] : 
                        (N179)? \xnz.mem_r [123] : 
                        (N181)? \xnz.mem_r [156] : 
                        (N183)? \xnz.mem_r [189] : 
                        (N185)? \xnz.mem_r [222] : 
                        (N187)? \xnz.mem_r [255] : 
                        (N189)? \xnz.mem_r [288] : 
                        (N191)? \xnz.mem_r [321] : 
                        (N193)? \xnz.mem_r [354] : 
                        (N195)? \xnz.mem_r [387] : 
                        (N197)? \xnz.mem_r [420] : 
                        (N199)? \xnz.mem_r [453] : 
                        (N201)? \xnz.mem_r [486] : 
                        (N203)? \xnz.mem_r [519] : 
                        (N174)? \xnz.mem_r [552] : 
                        (N176)? \xnz.mem_r [585] : 
                        (N178)? \xnz.mem_r [618] : 
                        (N180)? \xnz.mem_r [651] : 
                        (N182)? \xnz.mem_r [684] : 
                        (N184)? \xnz.mem_r [717] : 
                        (N186)? \xnz.mem_r [750] : 
                        (N188)? \xnz.mem_r [783] : 
                        (N190)? \xnz.mem_r [816] : 
                        (N192)? \xnz.mem_r [849] : 
                        (N194)? \xnz.mem_r [882] : 
                        (N196)? \xnz.mem_r [915] : 
                        (N198)? \xnz.mem_r [948] : 
                        (N200)? \xnz.mem_r [981] : 
                        (N202)? \xnz.mem_r [1014] : 
                        (N204)? \xnz.mem_r [1047] : 1'b0;
  assign r_data_o[89] = (N173)? \xnz.mem_r [23] : 
                        (N175)? \xnz.mem_r [56] : 
                        (N177)? \xnz.mem_r [89] : 
                        (N179)? \xnz.mem_r [122] : 
                        (N181)? \xnz.mem_r [155] : 
                        (N183)? \xnz.mem_r [188] : 
                        (N185)? \xnz.mem_r [221] : 
                        (N187)? \xnz.mem_r [254] : 
                        (N189)? \xnz.mem_r [287] : 
                        (N191)? \xnz.mem_r [320] : 
                        (N193)? \xnz.mem_r [353] : 
                        (N195)? \xnz.mem_r [386] : 
                        (N197)? \xnz.mem_r [419] : 
                        (N199)? \xnz.mem_r [452] : 
                        (N201)? \xnz.mem_r [485] : 
                        (N203)? \xnz.mem_r [518] : 
                        (N174)? \xnz.mem_r [551] : 
                        (N176)? \xnz.mem_r [584] : 
                        (N178)? \xnz.mem_r [617] : 
                        (N180)? \xnz.mem_r [650] : 
                        (N182)? \xnz.mem_r [683] : 
                        (N184)? \xnz.mem_r [716] : 
                        (N186)? \xnz.mem_r [749] : 
                        (N188)? \xnz.mem_r [782] : 
                        (N190)? \xnz.mem_r [815] : 
                        (N192)? \xnz.mem_r [848] : 
                        (N194)? \xnz.mem_r [881] : 
                        (N196)? \xnz.mem_r [914] : 
                        (N198)? \xnz.mem_r [947] : 
                        (N200)? \xnz.mem_r [980] : 
                        (N202)? \xnz.mem_r [1013] : 
                        (N204)? \xnz.mem_r [1046] : 1'b0;
  assign r_data_o[88] = (N173)? \xnz.mem_r [22] : 
                        (N175)? \xnz.mem_r [55] : 
                        (N177)? \xnz.mem_r [88] : 
                        (N179)? \xnz.mem_r [121] : 
                        (N181)? \xnz.mem_r [154] : 
                        (N183)? \xnz.mem_r [187] : 
                        (N185)? \xnz.mem_r [220] : 
                        (N187)? \xnz.mem_r [253] : 
                        (N189)? \xnz.mem_r [286] : 
                        (N191)? \xnz.mem_r [319] : 
                        (N193)? \xnz.mem_r [352] : 
                        (N195)? \xnz.mem_r [385] : 
                        (N197)? \xnz.mem_r [418] : 
                        (N199)? \xnz.mem_r [451] : 
                        (N201)? \xnz.mem_r [484] : 
                        (N203)? \xnz.mem_r [517] : 
                        (N174)? \xnz.mem_r [550] : 
                        (N176)? \xnz.mem_r [583] : 
                        (N178)? \xnz.mem_r [616] : 
                        (N180)? \xnz.mem_r [649] : 
                        (N182)? \xnz.mem_r [682] : 
                        (N184)? \xnz.mem_r [715] : 
                        (N186)? \xnz.mem_r [748] : 
                        (N188)? \xnz.mem_r [781] : 
                        (N190)? \xnz.mem_r [814] : 
                        (N192)? \xnz.mem_r [847] : 
                        (N194)? \xnz.mem_r [880] : 
                        (N196)? \xnz.mem_r [913] : 
                        (N198)? \xnz.mem_r [946] : 
                        (N200)? \xnz.mem_r [979] : 
                        (N202)? \xnz.mem_r [1012] : 
                        (N204)? \xnz.mem_r [1045] : 1'b0;
  assign r_data_o[87] = (N173)? \xnz.mem_r [21] : 
                        (N175)? \xnz.mem_r [54] : 
                        (N177)? \xnz.mem_r [87] : 
                        (N179)? \xnz.mem_r [120] : 
                        (N181)? \xnz.mem_r [153] : 
                        (N183)? \xnz.mem_r [186] : 
                        (N185)? \xnz.mem_r [219] : 
                        (N187)? \xnz.mem_r [252] : 
                        (N189)? \xnz.mem_r [285] : 
                        (N191)? \xnz.mem_r [318] : 
                        (N193)? \xnz.mem_r [351] : 
                        (N195)? \xnz.mem_r [384] : 
                        (N197)? \xnz.mem_r [417] : 
                        (N199)? \xnz.mem_r [450] : 
                        (N201)? \xnz.mem_r [483] : 
                        (N203)? \xnz.mem_r [516] : 
                        (N174)? \xnz.mem_r [549] : 
                        (N176)? \xnz.mem_r [582] : 
                        (N178)? \xnz.mem_r [615] : 
                        (N180)? \xnz.mem_r [648] : 
                        (N182)? \xnz.mem_r [681] : 
                        (N184)? \xnz.mem_r [714] : 
                        (N186)? \xnz.mem_r [747] : 
                        (N188)? \xnz.mem_r [780] : 
                        (N190)? \xnz.mem_r [813] : 
                        (N192)? \xnz.mem_r [846] : 
                        (N194)? \xnz.mem_r [879] : 
                        (N196)? \xnz.mem_r [912] : 
                        (N198)? \xnz.mem_r [945] : 
                        (N200)? \xnz.mem_r [978] : 
                        (N202)? \xnz.mem_r [1011] : 
                        (N204)? \xnz.mem_r [1044] : 1'b0;
  assign r_data_o[86] = (N173)? \xnz.mem_r [20] : 
                        (N175)? \xnz.mem_r [53] : 
                        (N177)? \xnz.mem_r [86] : 
                        (N179)? \xnz.mem_r [119] : 
                        (N181)? \xnz.mem_r [152] : 
                        (N183)? \xnz.mem_r [185] : 
                        (N185)? \xnz.mem_r [218] : 
                        (N187)? \xnz.mem_r [251] : 
                        (N189)? \xnz.mem_r [284] : 
                        (N191)? \xnz.mem_r [317] : 
                        (N193)? \xnz.mem_r [350] : 
                        (N195)? \xnz.mem_r [383] : 
                        (N197)? \xnz.mem_r [416] : 
                        (N199)? \xnz.mem_r [449] : 
                        (N201)? \xnz.mem_r [482] : 
                        (N203)? \xnz.mem_r [515] : 
                        (N174)? \xnz.mem_r [548] : 
                        (N176)? \xnz.mem_r [581] : 
                        (N178)? \xnz.mem_r [614] : 
                        (N180)? \xnz.mem_r [647] : 
                        (N182)? \xnz.mem_r [680] : 
                        (N184)? \xnz.mem_r [713] : 
                        (N186)? \xnz.mem_r [746] : 
                        (N188)? \xnz.mem_r [779] : 
                        (N190)? \xnz.mem_r [812] : 
                        (N192)? \xnz.mem_r [845] : 
                        (N194)? \xnz.mem_r [878] : 
                        (N196)? \xnz.mem_r [911] : 
                        (N198)? \xnz.mem_r [944] : 
                        (N200)? \xnz.mem_r [977] : 
                        (N202)? \xnz.mem_r [1010] : 
                        (N204)? \xnz.mem_r [1043] : 1'b0;
  assign r_data_o[85] = (N173)? \xnz.mem_r [19] : 
                        (N175)? \xnz.mem_r [52] : 
                        (N177)? \xnz.mem_r [85] : 
                        (N179)? \xnz.mem_r [118] : 
                        (N181)? \xnz.mem_r [151] : 
                        (N183)? \xnz.mem_r [184] : 
                        (N185)? \xnz.mem_r [217] : 
                        (N187)? \xnz.mem_r [250] : 
                        (N189)? \xnz.mem_r [283] : 
                        (N191)? \xnz.mem_r [316] : 
                        (N193)? \xnz.mem_r [349] : 
                        (N195)? \xnz.mem_r [382] : 
                        (N197)? \xnz.mem_r [415] : 
                        (N199)? \xnz.mem_r [448] : 
                        (N201)? \xnz.mem_r [481] : 
                        (N203)? \xnz.mem_r [514] : 
                        (N174)? \xnz.mem_r [547] : 
                        (N176)? \xnz.mem_r [580] : 
                        (N178)? \xnz.mem_r [613] : 
                        (N180)? \xnz.mem_r [646] : 
                        (N182)? \xnz.mem_r [679] : 
                        (N184)? \xnz.mem_r [712] : 
                        (N186)? \xnz.mem_r [745] : 
                        (N188)? \xnz.mem_r [778] : 
                        (N190)? \xnz.mem_r [811] : 
                        (N192)? \xnz.mem_r [844] : 
                        (N194)? \xnz.mem_r [877] : 
                        (N196)? \xnz.mem_r [910] : 
                        (N198)? \xnz.mem_r [943] : 
                        (N200)? \xnz.mem_r [976] : 
                        (N202)? \xnz.mem_r [1009] : 
                        (N204)? \xnz.mem_r [1042] : 1'b0;
  assign r_data_o[84] = (N173)? \xnz.mem_r [18] : 
                        (N175)? \xnz.mem_r [51] : 
                        (N177)? \xnz.mem_r [84] : 
                        (N179)? \xnz.mem_r [117] : 
                        (N181)? \xnz.mem_r [150] : 
                        (N183)? \xnz.mem_r [183] : 
                        (N185)? \xnz.mem_r [216] : 
                        (N187)? \xnz.mem_r [249] : 
                        (N189)? \xnz.mem_r [282] : 
                        (N191)? \xnz.mem_r [315] : 
                        (N193)? \xnz.mem_r [348] : 
                        (N195)? \xnz.mem_r [381] : 
                        (N197)? \xnz.mem_r [414] : 
                        (N199)? \xnz.mem_r [447] : 
                        (N201)? \xnz.mem_r [480] : 
                        (N203)? \xnz.mem_r [513] : 
                        (N174)? \xnz.mem_r [546] : 
                        (N176)? \xnz.mem_r [579] : 
                        (N178)? \xnz.mem_r [612] : 
                        (N180)? \xnz.mem_r [645] : 
                        (N182)? \xnz.mem_r [678] : 
                        (N184)? \xnz.mem_r [711] : 
                        (N186)? \xnz.mem_r [744] : 
                        (N188)? \xnz.mem_r [777] : 
                        (N190)? \xnz.mem_r [810] : 
                        (N192)? \xnz.mem_r [843] : 
                        (N194)? \xnz.mem_r [876] : 
                        (N196)? \xnz.mem_r [909] : 
                        (N198)? \xnz.mem_r [942] : 
                        (N200)? \xnz.mem_r [975] : 
                        (N202)? \xnz.mem_r [1008] : 
                        (N204)? \xnz.mem_r [1041] : 1'b0;
  assign r_data_o[83] = (N173)? \xnz.mem_r [17] : 
                        (N175)? \xnz.mem_r [50] : 
                        (N177)? \xnz.mem_r [83] : 
                        (N179)? \xnz.mem_r [116] : 
                        (N181)? \xnz.mem_r [149] : 
                        (N183)? \xnz.mem_r [182] : 
                        (N185)? \xnz.mem_r [215] : 
                        (N187)? \xnz.mem_r [248] : 
                        (N189)? \xnz.mem_r [281] : 
                        (N191)? \xnz.mem_r [314] : 
                        (N193)? \xnz.mem_r [347] : 
                        (N195)? \xnz.mem_r [380] : 
                        (N197)? \xnz.mem_r [413] : 
                        (N199)? \xnz.mem_r [446] : 
                        (N201)? \xnz.mem_r [479] : 
                        (N203)? \xnz.mem_r [512] : 
                        (N174)? \xnz.mem_r [545] : 
                        (N176)? \xnz.mem_r [578] : 
                        (N178)? \xnz.mem_r [611] : 
                        (N180)? \xnz.mem_r [644] : 
                        (N182)? \xnz.mem_r [677] : 
                        (N184)? \xnz.mem_r [710] : 
                        (N186)? \xnz.mem_r [743] : 
                        (N188)? \xnz.mem_r [776] : 
                        (N190)? \xnz.mem_r [809] : 
                        (N192)? \xnz.mem_r [842] : 
                        (N194)? \xnz.mem_r [875] : 
                        (N196)? \xnz.mem_r [908] : 
                        (N198)? \xnz.mem_r [941] : 
                        (N200)? \xnz.mem_r [974] : 
                        (N202)? \xnz.mem_r [1007] : 
                        (N204)? \xnz.mem_r [1040] : 1'b0;
  assign r_data_o[82] = (N173)? \xnz.mem_r [16] : 
                        (N175)? \xnz.mem_r [49] : 
                        (N177)? \xnz.mem_r [82] : 
                        (N179)? \xnz.mem_r [115] : 
                        (N181)? \xnz.mem_r [148] : 
                        (N183)? \xnz.mem_r [181] : 
                        (N185)? \xnz.mem_r [214] : 
                        (N187)? \xnz.mem_r [247] : 
                        (N189)? \xnz.mem_r [280] : 
                        (N191)? \xnz.mem_r [313] : 
                        (N193)? \xnz.mem_r [346] : 
                        (N195)? \xnz.mem_r [379] : 
                        (N197)? \xnz.mem_r [412] : 
                        (N199)? \xnz.mem_r [445] : 
                        (N201)? \xnz.mem_r [478] : 
                        (N203)? \xnz.mem_r [511] : 
                        (N174)? \xnz.mem_r [544] : 
                        (N176)? \xnz.mem_r [577] : 
                        (N178)? \xnz.mem_r [610] : 
                        (N180)? \xnz.mem_r [643] : 
                        (N182)? \xnz.mem_r [676] : 
                        (N184)? \xnz.mem_r [709] : 
                        (N186)? \xnz.mem_r [742] : 
                        (N188)? \xnz.mem_r [775] : 
                        (N190)? \xnz.mem_r [808] : 
                        (N192)? \xnz.mem_r [841] : 
                        (N194)? \xnz.mem_r [874] : 
                        (N196)? \xnz.mem_r [907] : 
                        (N198)? \xnz.mem_r [940] : 
                        (N200)? \xnz.mem_r [973] : 
                        (N202)? \xnz.mem_r [1006] : 
                        (N204)? \xnz.mem_r [1039] : 1'b0;
  assign r_data_o[81] = (N173)? \xnz.mem_r [15] : 
                        (N175)? \xnz.mem_r [48] : 
                        (N177)? \xnz.mem_r [81] : 
                        (N179)? \xnz.mem_r [114] : 
                        (N181)? \xnz.mem_r [147] : 
                        (N183)? \xnz.mem_r [180] : 
                        (N185)? \xnz.mem_r [213] : 
                        (N187)? \xnz.mem_r [246] : 
                        (N189)? \xnz.mem_r [279] : 
                        (N191)? \xnz.mem_r [312] : 
                        (N193)? \xnz.mem_r [345] : 
                        (N195)? \xnz.mem_r [378] : 
                        (N197)? \xnz.mem_r [411] : 
                        (N199)? \xnz.mem_r [444] : 
                        (N201)? \xnz.mem_r [477] : 
                        (N203)? \xnz.mem_r [510] : 
                        (N174)? \xnz.mem_r [543] : 
                        (N176)? \xnz.mem_r [576] : 
                        (N178)? \xnz.mem_r [609] : 
                        (N180)? \xnz.mem_r [642] : 
                        (N182)? \xnz.mem_r [675] : 
                        (N184)? \xnz.mem_r [708] : 
                        (N186)? \xnz.mem_r [741] : 
                        (N188)? \xnz.mem_r [774] : 
                        (N190)? \xnz.mem_r [807] : 
                        (N192)? \xnz.mem_r [840] : 
                        (N194)? \xnz.mem_r [873] : 
                        (N196)? \xnz.mem_r [906] : 
                        (N198)? \xnz.mem_r [939] : 
                        (N200)? \xnz.mem_r [972] : 
                        (N202)? \xnz.mem_r [1005] : 
                        (N204)? \xnz.mem_r [1038] : 1'b0;
  assign r_data_o[80] = (N173)? \xnz.mem_r [14] : 
                        (N175)? \xnz.mem_r [47] : 
                        (N177)? \xnz.mem_r [80] : 
                        (N179)? \xnz.mem_r [113] : 
                        (N181)? \xnz.mem_r [146] : 
                        (N183)? \xnz.mem_r [179] : 
                        (N185)? \xnz.mem_r [212] : 
                        (N187)? \xnz.mem_r [245] : 
                        (N189)? \xnz.mem_r [278] : 
                        (N191)? \xnz.mem_r [311] : 
                        (N193)? \xnz.mem_r [344] : 
                        (N195)? \xnz.mem_r [377] : 
                        (N197)? \xnz.mem_r [410] : 
                        (N199)? \xnz.mem_r [443] : 
                        (N201)? \xnz.mem_r [476] : 
                        (N203)? \xnz.mem_r [509] : 
                        (N174)? \xnz.mem_r [542] : 
                        (N176)? \xnz.mem_r [575] : 
                        (N178)? \xnz.mem_r [608] : 
                        (N180)? \xnz.mem_r [641] : 
                        (N182)? \xnz.mem_r [674] : 
                        (N184)? \xnz.mem_r [707] : 
                        (N186)? \xnz.mem_r [740] : 
                        (N188)? \xnz.mem_r [773] : 
                        (N190)? \xnz.mem_r [806] : 
                        (N192)? \xnz.mem_r [839] : 
                        (N194)? \xnz.mem_r [872] : 
                        (N196)? \xnz.mem_r [905] : 
                        (N198)? \xnz.mem_r [938] : 
                        (N200)? \xnz.mem_r [971] : 
                        (N202)? \xnz.mem_r [1004] : 
                        (N204)? \xnz.mem_r [1037] : 1'b0;
  assign r_data_o[79] = (N173)? \xnz.mem_r [13] : 
                        (N175)? \xnz.mem_r [46] : 
                        (N177)? \xnz.mem_r [79] : 
                        (N179)? \xnz.mem_r [112] : 
                        (N181)? \xnz.mem_r [145] : 
                        (N183)? \xnz.mem_r [178] : 
                        (N185)? \xnz.mem_r [211] : 
                        (N187)? \xnz.mem_r [244] : 
                        (N189)? \xnz.mem_r [277] : 
                        (N191)? \xnz.mem_r [310] : 
                        (N193)? \xnz.mem_r [343] : 
                        (N195)? \xnz.mem_r [376] : 
                        (N197)? \xnz.mem_r [409] : 
                        (N199)? \xnz.mem_r [442] : 
                        (N201)? \xnz.mem_r [475] : 
                        (N203)? \xnz.mem_r [508] : 
                        (N174)? \xnz.mem_r [541] : 
                        (N176)? \xnz.mem_r [574] : 
                        (N178)? \xnz.mem_r [607] : 
                        (N180)? \xnz.mem_r [640] : 
                        (N182)? \xnz.mem_r [673] : 
                        (N184)? \xnz.mem_r [706] : 
                        (N186)? \xnz.mem_r [739] : 
                        (N188)? \xnz.mem_r [772] : 
                        (N190)? \xnz.mem_r [805] : 
                        (N192)? \xnz.mem_r [838] : 
                        (N194)? \xnz.mem_r [871] : 
                        (N196)? \xnz.mem_r [904] : 
                        (N198)? \xnz.mem_r [937] : 
                        (N200)? \xnz.mem_r [970] : 
                        (N202)? \xnz.mem_r [1003] : 
                        (N204)? \xnz.mem_r [1036] : 1'b0;
  assign r_data_o[78] = (N173)? \xnz.mem_r [12] : 
                        (N175)? \xnz.mem_r [45] : 
                        (N177)? \xnz.mem_r [78] : 
                        (N179)? \xnz.mem_r [111] : 
                        (N181)? \xnz.mem_r [144] : 
                        (N183)? \xnz.mem_r [177] : 
                        (N185)? \xnz.mem_r [210] : 
                        (N187)? \xnz.mem_r [243] : 
                        (N189)? \xnz.mem_r [276] : 
                        (N191)? \xnz.mem_r [309] : 
                        (N193)? \xnz.mem_r [342] : 
                        (N195)? \xnz.mem_r [375] : 
                        (N197)? \xnz.mem_r [408] : 
                        (N199)? \xnz.mem_r [441] : 
                        (N201)? \xnz.mem_r [474] : 
                        (N203)? \xnz.mem_r [507] : 
                        (N174)? \xnz.mem_r [540] : 
                        (N176)? \xnz.mem_r [573] : 
                        (N178)? \xnz.mem_r [606] : 
                        (N180)? \xnz.mem_r [639] : 
                        (N182)? \xnz.mem_r [672] : 
                        (N184)? \xnz.mem_r [705] : 
                        (N186)? \xnz.mem_r [738] : 
                        (N188)? \xnz.mem_r [771] : 
                        (N190)? \xnz.mem_r [804] : 
                        (N192)? \xnz.mem_r [837] : 
                        (N194)? \xnz.mem_r [870] : 
                        (N196)? \xnz.mem_r [903] : 
                        (N198)? \xnz.mem_r [936] : 
                        (N200)? \xnz.mem_r [969] : 
                        (N202)? \xnz.mem_r [1002] : 
                        (N204)? \xnz.mem_r [1035] : 1'b0;
  assign r_data_o[77] = (N173)? \xnz.mem_r [11] : 
                        (N175)? \xnz.mem_r [44] : 
                        (N177)? \xnz.mem_r [77] : 
                        (N179)? \xnz.mem_r [110] : 
                        (N181)? \xnz.mem_r [143] : 
                        (N183)? \xnz.mem_r [176] : 
                        (N185)? \xnz.mem_r [209] : 
                        (N187)? \xnz.mem_r [242] : 
                        (N189)? \xnz.mem_r [275] : 
                        (N191)? \xnz.mem_r [308] : 
                        (N193)? \xnz.mem_r [341] : 
                        (N195)? \xnz.mem_r [374] : 
                        (N197)? \xnz.mem_r [407] : 
                        (N199)? \xnz.mem_r [440] : 
                        (N201)? \xnz.mem_r [473] : 
                        (N203)? \xnz.mem_r [506] : 
                        (N174)? \xnz.mem_r [539] : 
                        (N176)? \xnz.mem_r [572] : 
                        (N178)? \xnz.mem_r [605] : 
                        (N180)? \xnz.mem_r [638] : 
                        (N182)? \xnz.mem_r [671] : 
                        (N184)? \xnz.mem_r [704] : 
                        (N186)? \xnz.mem_r [737] : 
                        (N188)? \xnz.mem_r [770] : 
                        (N190)? \xnz.mem_r [803] : 
                        (N192)? \xnz.mem_r [836] : 
                        (N194)? \xnz.mem_r [869] : 
                        (N196)? \xnz.mem_r [902] : 
                        (N198)? \xnz.mem_r [935] : 
                        (N200)? \xnz.mem_r [968] : 
                        (N202)? \xnz.mem_r [1001] : 
                        (N204)? \xnz.mem_r [1034] : 1'b0;
  assign r_data_o[76] = (N173)? \xnz.mem_r [10] : 
                        (N175)? \xnz.mem_r [43] : 
                        (N177)? \xnz.mem_r [76] : 
                        (N179)? \xnz.mem_r [109] : 
                        (N181)? \xnz.mem_r [142] : 
                        (N183)? \xnz.mem_r [175] : 
                        (N185)? \xnz.mem_r [208] : 
                        (N187)? \xnz.mem_r [241] : 
                        (N189)? \xnz.mem_r [274] : 
                        (N191)? \xnz.mem_r [307] : 
                        (N193)? \xnz.mem_r [340] : 
                        (N195)? \xnz.mem_r [373] : 
                        (N197)? \xnz.mem_r [406] : 
                        (N199)? \xnz.mem_r [439] : 
                        (N201)? \xnz.mem_r [472] : 
                        (N203)? \xnz.mem_r [505] : 
                        (N174)? \xnz.mem_r [538] : 
                        (N176)? \xnz.mem_r [571] : 
                        (N178)? \xnz.mem_r [604] : 
                        (N180)? \xnz.mem_r [637] : 
                        (N182)? \xnz.mem_r [670] : 
                        (N184)? \xnz.mem_r [703] : 
                        (N186)? \xnz.mem_r [736] : 
                        (N188)? \xnz.mem_r [769] : 
                        (N190)? \xnz.mem_r [802] : 
                        (N192)? \xnz.mem_r [835] : 
                        (N194)? \xnz.mem_r [868] : 
                        (N196)? \xnz.mem_r [901] : 
                        (N198)? \xnz.mem_r [934] : 
                        (N200)? \xnz.mem_r [967] : 
                        (N202)? \xnz.mem_r [1000] : 
                        (N204)? \xnz.mem_r [1033] : 1'b0;
  assign r_data_o[75] = (N173)? \xnz.mem_r [9] : 
                        (N175)? \xnz.mem_r [42] : 
                        (N177)? \xnz.mem_r [75] : 
                        (N179)? \xnz.mem_r [108] : 
                        (N181)? \xnz.mem_r [141] : 
                        (N183)? \xnz.mem_r [174] : 
                        (N185)? \xnz.mem_r [207] : 
                        (N187)? \xnz.mem_r [240] : 
                        (N189)? \xnz.mem_r [273] : 
                        (N191)? \xnz.mem_r [306] : 
                        (N193)? \xnz.mem_r [339] : 
                        (N195)? \xnz.mem_r [372] : 
                        (N197)? \xnz.mem_r [405] : 
                        (N199)? \xnz.mem_r [438] : 
                        (N201)? \xnz.mem_r [471] : 
                        (N203)? \xnz.mem_r [504] : 
                        (N174)? \xnz.mem_r [537] : 
                        (N176)? \xnz.mem_r [570] : 
                        (N178)? \xnz.mem_r [603] : 
                        (N180)? \xnz.mem_r [636] : 
                        (N182)? \xnz.mem_r [669] : 
                        (N184)? \xnz.mem_r [702] : 
                        (N186)? \xnz.mem_r [735] : 
                        (N188)? \xnz.mem_r [768] : 
                        (N190)? \xnz.mem_r [801] : 
                        (N192)? \xnz.mem_r [834] : 
                        (N194)? \xnz.mem_r [867] : 
                        (N196)? \xnz.mem_r [900] : 
                        (N198)? \xnz.mem_r [933] : 
                        (N200)? \xnz.mem_r [966] : 
                        (N202)? \xnz.mem_r [999] : 
                        (N204)? \xnz.mem_r [1032] : 1'b0;
  assign r_data_o[74] = (N173)? \xnz.mem_r [8] : 
                        (N175)? \xnz.mem_r [41] : 
                        (N177)? \xnz.mem_r [74] : 
                        (N179)? \xnz.mem_r [107] : 
                        (N181)? \xnz.mem_r [140] : 
                        (N183)? \xnz.mem_r [173] : 
                        (N185)? \xnz.mem_r [206] : 
                        (N187)? \xnz.mem_r [239] : 
                        (N189)? \xnz.mem_r [272] : 
                        (N191)? \xnz.mem_r [305] : 
                        (N193)? \xnz.mem_r [338] : 
                        (N195)? \xnz.mem_r [371] : 
                        (N197)? \xnz.mem_r [404] : 
                        (N199)? \xnz.mem_r [437] : 
                        (N201)? \xnz.mem_r [470] : 
                        (N203)? \xnz.mem_r [503] : 
                        (N174)? \xnz.mem_r [536] : 
                        (N176)? \xnz.mem_r [569] : 
                        (N178)? \xnz.mem_r [602] : 
                        (N180)? \xnz.mem_r [635] : 
                        (N182)? \xnz.mem_r [668] : 
                        (N184)? \xnz.mem_r [701] : 
                        (N186)? \xnz.mem_r [734] : 
                        (N188)? \xnz.mem_r [767] : 
                        (N190)? \xnz.mem_r [800] : 
                        (N192)? \xnz.mem_r [833] : 
                        (N194)? \xnz.mem_r [866] : 
                        (N196)? \xnz.mem_r [899] : 
                        (N198)? \xnz.mem_r [932] : 
                        (N200)? \xnz.mem_r [965] : 
                        (N202)? \xnz.mem_r [998] : 
                        (N204)? \xnz.mem_r [1031] : 1'b0;
  assign r_data_o[73] = (N173)? \xnz.mem_r [7] : 
                        (N175)? \xnz.mem_r [40] : 
                        (N177)? \xnz.mem_r [73] : 
                        (N179)? \xnz.mem_r [106] : 
                        (N181)? \xnz.mem_r [139] : 
                        (N183)? \xnz.mem_r [172] : 
                        (N185)? \xnz.mem_r [205] : 
                        (N187)? \xnz.mem_r [238] : 
                        (N189)? \xnz.mem_r [271] : 
                        (N191)? \xnz.mem_r [304] : 
                        (N193)? \xnz.mem_r [337] : 
                        (N195)? \xnz.mem_r [370] : 
                        (N197)? \xnz.mem_r [403] : 
                        (N199)? \xnz.mem_r [436] : 
                        (N201)? \xnz.mem_r [469] : 
                        (N203)? \xnz.mem_r [502] : 
                        (N174)? \xnz.mem_r [535] : 
                        (N176)? \xnz.mem_r [568] : 
                        (N178)? \xnz.mem_r [601] : 
                        (N180)? \xnz.mem_r [634] : 
                        (N182)? \xnz.mem_r [667] : 
                        (N184)? \xnz.mem_r [700] : 
                        (N186)? \xnz.mem_r [733] : 
                        (N188)? \xnz.mem_r [766] : 
                        (N190)? \xnz.mem_r [799] : 
                        (N192)? \xnz.mem_r [832] : 
                        (N194)? \xnz.mem_r [865] : 
                        (N196)? \xnz.mem_r [898] : 
                        (N198)? \xnz.mem_r [931] : 
                        (N200)? \xnz.mem_r [964] : 
                        (N202)? \xnz.mem_r [997] : 
                        (N204)? \xnz.mem_r [1030] : 1'b0;
  assign r_data_o[72] = (N173)? \xnz.mem_r [6] : 
                        (N175)? \xnz.mem_r [39] : 
                        (N177)? \xnz.mem_r [72] : 
                        (N179)? \xnz.mem_r [105] : 
                        (N181)? \xnz.mem_r [138] : 
                        (N183)? \xnz.mem_r [171] : 
                        (N185)? \xnz.mem_r [204] : 
                        (N187)? \xnz.mem_r [237] : 
                        (N189)? \xnz.mem_r [270] : 
                        (N191)? \xnz.mem_r [303] : 
                        (N193)? \xnz.mem_r [336] : 
                        (N195)? \xnz.mem_r [369] : 
                        (N197)? \xnz.mem_r [402] : 
                        (N199)? \xnz.mem_r [435] : 
                        (N201)? \xnz.mem_r [468] : 
                        (N203)? \xnz.mem_r [501] : 
                        (N174)? \xnz.mem_r [534] : 
                        (N176)? \xnz.mem_r [567] : 
                        (N178)? \xnz.mem_r [600] : 
                        (N180)? \xnz.mem_r [633] : 
                        (N182)? \xnz.mem_r [666] : 
                        (N184)? \xnz.mem_r [699] : 
                        (N186)? \xnz.mem_r [732] : 
                        (N188)? \xnz.mem_r [765] : 
                        (N190)? \xnz.mem_r [798] : 
                        (N192)? \xnz.mem_r [831] : 
                        (N194)? \xnz.mem_r [864] : 
                        (N196)? \xnz.mem_r [897] : 
                        (N198)? \xnz.mem_r [930] : 
                        (N200)? \xnz.mem_r [963] : 
                        (N202)? \xnz.mem_r [996] : 
                        (N204)? \xnz.mem_r [1029] : 1'b0;
  assign r_data_o[71] = (N173)? \xnz.mem_r [5] : 
                        (N175)? \xnz.mem_r [38] : 
                        (N177)? \xnz.mem_r [71] : 
                        (N179)? \xnz.mem_r [104] : 
                        (N181)? \xnz.mem_r [137] : 
                        (N183)? \xnz.mem_r [170] : 
                        (N185)? \xnz.mem_r [203] : 
                        (N187)? \xnz.mem_r [236] : 
                        (N189)? \xnz.mem_r [269] : 
                        (N191)? \xnz.mem_r [302] : 
                        (N193)? \xnz.mem_r [335] : 
                        (N195)? \xnz.mem_r [368] : 
                        (N197)? \xnz.mem_r [401] : 
                        (N199)? \xnz.mem_r [434] : 
                        (N201)? \xnz.mem_r [467] : 
                        (N203)? \xnz.mem_r [500] : 
                        (N174)? \xnz.mem_r [533] : 
                        (N176)? \xnz.mem_r [566] : 
                        (N178)? \xnz.mem_r [599] : 
                        (N180)? \xnz.mem_r [632] : 
                        (N182)? \xnz.mem_r [665] : 
                        (N184)? \xnz.mem_r [698] : 
                        (N186)? \xnz.mem_r [731] : 
                        (N188)? \xnz.mem_r [764] : 
                        (N190)? \xnz.mem_r [797] : 
                        (N192)? \xnz.mem_r [830] : 
                        (N194)? \xnz.mem_r [863] : 
                        (N196)? \xnz.mem_r [896] : 
                        (N198)? \xnz.mem_r [929] : 
                        (N200)? \xnz.mem_r [962] : 
                        (N202)? \xnz.mem_r [995] : 
                        (N204)? \xnz.mem_r [1028] : 1'b0;
  assign r_data_o[70] = (N173)? \xnz.mem_r [4] : 
                        (N175)? \xnz.mem_r [37] : 
                        (N177)? \xnz.mem_r [70] : 
                        (N179)? \xnz.mem_r [103] : 
                        (N181)? \xnz.mem_r [136] : 
                        (N183)? \xnz.mem_r [169] : 
                        (N185)? \xnz.mem_r [202] : 
                        (N187)? \xnz.mem_r [235] : 
                        (N189)? \xnz.mem_r [268] : 
                        (N191)? \xnz.mem_r [301] : 
                        (N193)? \xnz.mem_r [334] : 
                        (N195)? \xnz.mem_r [367] : 
                        (N197)? \xnz.mem_r [400] : 
                        (N199)? \xnz.mem_r [433] : 
                        (N201)? \xnz.mem_r [466] : 
                        (N203)? \xnz.mem_r [499] : 
                        (N174)? \xnz.mem_r [532] : 
                        (N176)? \xnz.mem_r [565] : 
                        (N178)? \xnz.mem_r [598] : 
                        (N180)? \xnz.mem_r [631] : 
                        (N182)? \xnz.mem_r [664] : 
                        (N184)? \xnz.mem_r [697] : 
                        (N186)? \xnz.mem_r [730] : 
                        (N188)? \xnz.mem_r [763] : 
                        (N190)? \xnz.mem_r [796] : 
                        (N192)? \xnz.mem_r [829] : 
                        (N194)? \xnz.mem_r [862] : 
                        (N196)? \xnz.mem_r [895] : 
                        (N198)? \xnz.mem_r [928] : 
                        (N200)? \xnz.mem_r [961] : 
                        (N202)? \xnz.mem_r [994] : 
                        (N204)? \xnz.mem_r [1027] : 1'b0;
  assign r_data_o[69] = (N173)? \xnz.mem_r [3] : 
                        (N175)? \xnz.mem_r [36] : 
                        (N177)? \xnz.mem_r [69] : 
                        (N179)? \xnz.mem_r [102] : 
                        (N181)? \xnz.mem_r [135] : 
                        (N183)? \xnz.mem_r [168] : 
                        (N185)? \xnz.mem_r [201] : 
                        (N187)? \xnz.mem_r [234] : 
                        (N189)? \xnz.mem_r [267] : 
                        (N191)? \xnz.mem_r [300] : 
                        (N193)? \xnz.mem_r [333] : 
                        (N195)? \xnz.mem_r [366] : 
                        (N197)? \xnz.mem_r [399] : 
                        (N199)? \xnz.mem_r [432] : 
                        (N201)? \xnz.mem_r [465] : 
                        (N203)? \xnz.mem_r [498] : 
                        (N174)? \xnz.mem_r [531] : 
                        (N176)? \xnz.mem_r [564] : 
                        (N178)? \xnz.mem_r [597] : 
                        (N180)? \xnz.mem_r [630] : 
                        (N182)? \xnz.mem_r [663] : 
                        (N184)? \xnz.mem_r [696] : 
                        (N186)? \xnz.mem_r [729] : 
                        (N188)? \xnz.mem_r [762] : 
                        (N190)? \xnz.mem_r [795] : 
                        (N192)? \xnz.mem_r [828] : 
                        (N194)? \xnz.mem_r [861] : 
                        (N196)? \xnz.mem_r [894] : 
                        (N198)? \xnz.mem_r [927] : 
                        (N200)? \xnz.mem_r [960] : 
                        (N202)? \xnz.mem_r [993] : 
                        (N204)? \xnz.mem_r [1026] : 1'b0;
  assign r_data_o[68] = (N173)? \xnz.mem_r [2] : 
                        (N175)? \xnz.mem_r [35] : 
                        (N177)? \xnz.mem_r [68] : 
                        (N179)? \xnz.mem_r [101] : 
                        (N181)? \xnz.mem_r [134] : 
                        (N183)? \xnz.mem_r [167] : 
                        (N185)? \xnz.mem_r [200] : 
                        (N187)? \xnz.mem_r [233] : 
                        (N189)? \xnz.mem_r [266] : 
                        (N191)? \xnz.mem_r [299] : 
                        (N193)? \xnz.mem_r [332] : 
                        (N195)? \xnz.mem_r [365] : 
                        (N197)? \xnz.mem_r [398] : 
                        (N199)? \xnz.mem_r [431] : 
                        (N201)? \xnz.mem_r [464] : 
                        (N203)? \xnz.mem_r [497] : 
                        (N174)? \xnz.mem_r [530] : 
                        (N176)? \xnz.mem_r [563] : 
                        (N178)? \xnz.mem_r [596] : 
                        (N180)? \xnz.mem_r [629] : 
                        (N182)? \xnz.mem_r [662] : 
                        (N184)? \xnz.mem_r [695] : 
                        (N186)? \xnz.mem_r [728] : 
                        (N188)? \xnz.mem_r [761] : 
                        (N190)? \xnz.mem_r [794] : 
                        (N192)? \xnz.mem_r [827] : 
                        (N194)? \xnz.mem_r [860] : 
                        (N196)? \xnz.mem_r [893] : 
                        (N198)? \xnz.mem_r [926] : 
                        (N200)? \xnz.mem_r [959] : 
                        (N202)? \xnz.mem_r [992] : 
                        (N204)? \xnz.mem_r [1025] : 1'b0;
  assign r_data_o[67] = (N173)? \xnz.mem_r [1] : 
                        (N175)? \xnz.mem_r [34] : 
                        (N177)? \xnz.mem_r [67] : 
                        (N179)? \xnz.mem_r [100] : 
                        (N181)? \xnz.mem_r [133] : 
                        (N183)? \xnz.mem_r [166] : 
                        (N185)? \xnz.mem_r [199] : 
                        (N187)? \xnz.mem_r [232] : 
                        (N189)? \xnz.mem_r [265] : 
                        (N191)? \xnz.mem_r [298] : 
                        (N193)? \xnz.mem_r [331] : 
                        (N195)? \xnz.mem_r [364] : 
                        (N197)? \xnz.mem_r [397] : 
                        (N199)? \xnz.mem_r [430] : 
                        (N201)? \xnz.mem_r [463] : 
                        (N203)? \xnz.mem_r [496] : 
                        (N174)? \xnz.mem_r [529] : 
                        (N176)? \xnz.mem_r [562] : 
                        (N178)? \xnz.mem_r [595] : 
                        (N180)? \xnz.mem_r [628] : 
                        (N182)? \xnz.mem_r [661] : 
                        (N184)? \xnz.mem_r [694] : 
                        (N186)? \xnz.mem_r [727] : 
                        (N188)? \xnz.mem_r [760] : 
                        (N190)? \xnz.mem_r [793] : 
                        (N192)? \xnz.mem_r [826] : 
                        (N194)? \xnz.mem_r [859] : 
                        (N196)? \xnz.mem_r [892] : 
                        (N198)? \xnz.mem_r [925] : 
                        (N200)? \xnz.mem_r [958] : 
                        (N202)? \xnz.mem_r [991] : 
                        (N204)? \xnz.mem_r [1024] : 1'b0;
  assign r_data_o[66] = (N173)? \xnz.mem_r [0] : 
                        (N175)? \xnz.mem_r [33] : 
                        (N177)? \xnz.mem_r [66] : 
                        (N179)? \xnz.mem_r [99] : 
                        (N181)? \xnz.mem_r [132] : 
                        (N183)? \xnz.mem_r [165] : 
                        (N185)? \xnz.mem_r [198] : 
                        (N187)? \xnz.mem_r [231] : 
                        (N189)? \xnz.mem_r [264] : 
                        (N191)? \xnz.mem_r [297] : 
                        (N193)? \xnz.mem_r [330] : 
                        (N195)? \xnz.mem_r [363] : 
                        (N197)? \xnz.mem_r [396] : 
                        (N199)? \xnz.mem_r [429] : 
                        (N201)? \xnz.mem_r [462] : 
                        (N203)? \xnz.mem_r [495] : 
                        (N174)? \xnz.mem_r [528] : 
                        (N176)? \xnz.mem_r [561] : 
                        (N178)? \xnz.mem_r [594] : 
                        (N180)? \xnz.mem_r [627] : 
                        (N182)? \xnz.mem_r [660] : 
                        (N184)? \xnz.mem_r [693] : 
                        (N186)? \xnz.mem_r [726] : 
                        (N188)? \xnz.mem_r [759] : 
                        (N190)? \xnz.mem_r [792] : 
                        (N192)? \xnz.mem_r [825] : 
                        (N194)? \xnz.mem_r [858] : 
                        (N196)? \xnz.mem_r [891] : 
                        (N198)? \xnz.mem_r [924] : 
                        (N200)? \xnz.mem_r [957] : 
                        (N202)? \xnz.mem_r [990] : 
                        (N204)? \xnz.mem_r [1023] : 1'b0;
  assign N270 = w_addr_i[3] & w_addr_i[4];
  assign N271 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N272 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N273 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N274 = ~w_addr_i[2];
  assign N275 = w_addr_i[0] & w_addr_i[1];
  assign N276 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N277 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N278 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N279 = w_addr_i[2] & N275;
  assign N280 = w_addr_i[2] & N276;
  assign N281 = w_addr_i[2] & N277;
  assign N282 = w_addr_i[2] & N278;
  assign N283 = N274 & N275;
  assign N284 = N274 & N276;
  assign N285 = N274 & N277;
  assign N286 = N274 & N278;
  assign N237 = N270 & N279;
  assign N236 = N270 & N280;
  assign N235 = N270 & N281;
  assign N234 = N270 & N282;
  assign N233 = N270 & N283;
  assign N232 = N270 & N284;
  assign N231 = N270 & N285;
  assign N230 = N270 & N286;
  assign N229 = N271 & N279;
  assign N228 = N271 & N280;
  assign N227 = N271 & N281;
  assign N226 = N271 & N282;
  assign N225 = N271 & N283;
  assign N224 = N271 & N284;
  assign N223 = N271 & N285;
  assign N222 = N271 & N286;
  assign N221 = N272 & N279;
  assign N220 = N272 & N280;
  assign N219 = N272 & N281;
  assign N218 = N272 & N282;
  assign N217 = N272 & N283;
  assign N216 = N272 & N284;
  assign N215 = N272 & N285;
  assign N214 = N272 & N286;
  assign N213 = N273 & N279;
  assign N212 = N273 & N280;
  assign N211 = N273 & N281;
  assign N210 = N273 & N282;
  assign N209 = N273 & N283;
  assign N208 = N273 & N284;
  assign N207 = N273 & N285;
  assign N206 = N273 & N286;
  assign { N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238 } = (N8)? { N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206 } : 
                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N205;
  assign N10 = ~r_addr_r[0];
  assign N11 = ~r_addr_r[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_r[1];
  assign N14 = r_addr_r[0] & N11;
  assign N15 = r_addr_r[0] & r_addr_r[1];
  assign N16 = ~r_addr_r[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_r[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_r[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_r[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_r[2];
  assign N25 = ~r_addr_r[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_r[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_r[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_r[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_r[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_r[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_r[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_r[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_r[3];
  assign N42 = ~r_addr_r[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r_addr_r[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r_addr_r[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r_addr_r[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r_addr_r[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r_addr_r[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r_addr_r[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r_addr_r[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r_addr_r[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r_addr_r[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r_addr_r[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r_addr_r[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r_addr_r[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r_addr_r[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r_addr_r[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r_addr_r[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r_addr_r[4];
  assign N75 = ~r_addr_r[5];
  assign N76 = ~r_addr_r[6];
  assign N77 = N75 & N76;
  assign N78 = N75 & r_addr_r[6];
  assign N79 = r_addr_r[5] & N76;
  assign N80 = r_addr_r[5] & r_addr_r[6];
  assign N81 = ~r_addr_r[7];
  assign N82 = N77 & N81;
  assign N83 = N77 & r_addr_r[7];
  assign N84 = N79 & N81;
  assign N85 = N79 & r_addr_r[7];
  assign N86 = N78 & N81;
  assign N87 = N78 & r_addr_r[7];
  assign N88 = N80 & N81;
  assign N89 = N80 & r_addr_r[7];
  assign N90 = ~r_addr_r[8];
  assign N91 = N82 & N90;
  assign N92 = N82 & r_addr_r[8];
  assign N93 = N84 & N90;
  assign N94 = N84 & r_addr_r[8];
  assign N95 = N86 & N90;
  assign N96 = N86 & r_addr_r[8];
  assign N97 = N88 & N90;
  assign N98 = N88 & r_addr_r[8];
  assign N99 = N83 & N90;
  assign N100 = N83 & r_addr_r[8];
  assign N101 = N85 & N90;
  assign N102 = N85 & r_addr_r[8];
  assign N103 = N87 & N90;
  assign N104 = N87 & r_addr_r[8];
  assign N105 = N89 & N90;
  assign N106 = N89 & r_addr_r[8];
  assign N107 = ~r_addr_r[9];
  assign N108 = N91 & N107;
  assign N109 = N91 & r_addr_r[9];
  assign N110 = N93 & N107;
  assign N111 = N93 & r_addr_r[9];
  assign N112 = N95 & N107;
  assign N113 = N95 & r_addr_r[9];
  assign N114 = N97 & N107;
  assign N115 = N97 & r_addr_r[9];
  assign N116 = N99 & N107;
  assign N117 = N99 & r_addr_r[9];
  assign N118 = N101 & N107;
  assign N119 = N101 & r_addr_r[9];
  assign N120 = N103 & N107;
  assign N121 = N103 & r_addr_r[9];
  assign N122 = N105 & N107;
  assign N123 = N105 & r_addr_r[9];
  assign N124 = N92 & N107;
  assign N125 = N92 & r_addr_r[9];
  assign N126 = N94 & N107;
  assign N127 = N94 & r_addr_r[9];
  assign N128 = N96 & N107;
  assign N129 = N96 & r_addr_r[9];
  assign N130 = N98 & N107;
  assign N131 = N98 & r_addr_r[9];
  assign N132 = N100 & N107;
  assign N133 = N100 & r_addr_r[9];
  assign N134 = N102 & N107;
  assign N135 = N102 & r_addr_r[9];
  assign N136 = N104 & N107;
  assign N137 = N104 & r_addr_r[9];
  assign N138 = N106 & N107;
  assign N139 = N106 & r_addr_r[9];
  assign N140 = ~r_addr_r[10];
  assign N141 = ~r_addr_r[11];
  assign N142 = N140 & N141;
  assign N143 = N140 & r_addr_r[11];
  assign N144 = r_addr_r[10] & N141;
  assign N145 = r_addr_r[10] & r_addr_r[11];
  assign N146 = ~r_addr_r[12];
  assign N147 = N142 & N146;
  assign N148 = N142 & r_addr_r[12];
  assign N149 = N144 & N146;
  assign N150 = N144 & r_addr_r[12];
  assign N151 = N143 & N146;
  assign N152 = N143 & r_addr_r[12];
  assign N153 = N145 & N146;
  assign N154 = N145 & r_addr_r[12];
  assign N155 = ~r_addr_r[13];
  assign N156 = N147 & N155;
  assign N157 = N147 & r_addr_r[13];
  assign N158 = N149 & N155;
  assign N159 = N149 & r_addr_r[13];
  assign N160 = N151 & N155;
  assign N161 = N151 & r_addr_r[13];
  assign N162 = N153 & N155;
  assign N163 = N153 & r_addr_r[13];
  assign N164 = N148 & N155;
  assign N165 = N148 & r_addr_r[13];
  assign N166 = N150 & N155;
  assign N167 = N150 & r_addr_r[13];
  assign N168 = N152 & N155;
  assign N169 = N152 & r_addr_r[13];
  assign N170 = N154 & N155;
  assign N171 = N154 & r_addr_r[13];
  assign N172 = ~r_addr_r[14];
  assign N173 = N156 & N172;
  assign N174 = N156 & r_addr_r[14];
  assign N175 = N158 & N172;
  assign N176 = N158 & r_addr_r[14];
  assign N177 = N160 & N172;
  assign N178 = N160 & r_addr_r[14];
  assign N179 = N162 & N172;
  assign N180 = N162 & r_addr_r[14];
  assign N181 = N164 & N172;
  assign N182 = N164 & r_addr_r[14];
  assign N183 = N166 & N172;
  assign N184 = N166 & r_addr_r[14];
  assign N185 = N168 & N172;
  assign N186 = N168 & r_addr_r[14];
  assign N187 = N170 & N172;
  assign N188 = N170 & r_addr_r[14];
  assign N189 = N157 & N172;
  assign N190 = N157 & r_addr_r[14];
  assign N191 = N159 & N172;
  assign N192 = N159 & r_addr_r[14];
  assign N193 = N161 & N172;
  assign N194 = N161 & r_addr_r[14];
  assign N195 = N163 & N172;
  assign N196 = N163 & r_addr_r[14];
  assign N197 = N165 & N172;
  assign N198 = N165 & r_addr_r[14];
  assign N199 = N167 & N172;
  assign N200 = N167 & r_addr_r[14];
  assign N201 = N169 & N172;
  assign N202 = N169 & r_addr_r[14];
  assign N203 = N171 & N172;
  assign N204 = N171 & r_addr_r[14];
  assign N205 = ~w_v_i;

  always @(posedge clk_i) begin
    if(r_v_i[2]) begin
      r_addr_r_14_sv2v_reg <= r_addr_i[14];
      r_addr_r_13_sv2v_reg <= r_addr_i[13];
      r_addr_r_12_sv2v_reg <= r_addr_i[12];
      r_addr_r_11_sv2v_reg <= r_addr_i[11];
      r_addr_r_10_sv2v_reg <= r_addr_i[10];
    end 
    if(r_v_i[1]) begin
      r_addr_r_9_sv2v_reg <= r_addr_i[9];
      r_addr_r_8_sv2v_reg <= r_addr_i[8];
      r_addr_r_7_sv2v_reg <= r_addr_i[7];
      r_addr_r_6_sv2v_reg <= r_addr_i[6];
      r_addr_r_5_sv2v_reg <= r_addr_i[5];
    end 
    if(r_v_i[0]) begin
      r_addr_r_4_sv2v_reg <= r_addr_i[4];
      r_addr_r_3_sv2v_reg <= r_addr_i[3];
      r_addr_r_2_sv2v_reg <= r_addr_i[2];
      r_addr_r_1_sv2v_reg <= r_addr_i[1];
      r_addr_r_0_sv2v_reg <= r_addr_i[0];
    end 
    if(N269) begin
      \xnz.mem_r_1055_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_1054_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_1053_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_1052_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_1051_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_1050_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_1049_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_1048_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_1047_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_1046_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_1045_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_1044_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_1043_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_1042_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_1041_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_1040_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_1039_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_1038_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_1037_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_1036_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_1035_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_1034_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_1033_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_1032_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_1031_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_1030_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_1029_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_1028_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_1027_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_1026_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_1025_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_1024_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_1023_sv2v_reg  <= w_data_i[0];
    end 
    if(N268) begin
      \xnz.mem_r_1022_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_1021_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_1020_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_1019_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_1018_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_1017_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_1016_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_1015_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_1014_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_1013_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_1012_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_1011_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_1010_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_1009_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_1008_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_1007_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_1006_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_1005_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_1004_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_1003_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_1002_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_1001_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_1000_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_999_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_998_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_997_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_996_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_995_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_994_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_993_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_992_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_991_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_990_sv2v_reg  <= w_data_i[0];
    end 
    if(N267) begin
      \xnz.mem_r_989_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_988_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_987_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_986_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_985_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_984_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_983_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_982_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_981_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_980_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_979_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_978_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_977_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_976_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_975_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_974_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_973_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_972_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_971_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_970_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_969_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_968_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_967_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_966_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_965_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_964_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_963_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_962_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_961_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_960_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_959_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_958_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_957_sv2v_reg  <= w_data_i[0];
    end 
    if(N266) begin
      \xnz.mem_r_956_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_955_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_954_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_953_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_952_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_951_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_950_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_949_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_948_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_947_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_946_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_945_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_944_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_943_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_942_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_941_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_940_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_939_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_938_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_937_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_936_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_935_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_934_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_933_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_932_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_931_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_930_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_929_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_928_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_927_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_926_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_925_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_924_sv2v_reg  <= w_data_i[0];
    end 
    if(N265) begin
      \xnz.mem_r_923_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_922_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_921_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_920_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_919_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_918_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_917_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_916_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_915_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_914_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_913_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_912_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_911_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_910_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_909_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_908_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_907_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_906_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_905_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_904_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_903_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_902_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_901_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_900_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_899_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_898_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_897_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_896_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_895_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_894_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_893_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_892_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_891_sv2v_reg  <= w_data_i[0];
    end 
    if(N264) begin
      \xnz.mem_r_890_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_889_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_888_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_887_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_886_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_885_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_884_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_883_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_882_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_881_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_880_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_879_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_878_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_877_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_876_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_875_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_874_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_873_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_872_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_871_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_870_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_869_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_868_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_867_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_866_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_865_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_864_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_863_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_862_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_861_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_860_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_859_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_858_sv2v_reg  <= w_data_i[0];
    end 
    if(N263) begin
      \xnz.mem_r_857_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_856_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_855_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_854_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_853_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_852_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_851_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_850_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_849_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_848_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_847_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_846_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_845_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_844_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_843_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_842_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_841_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_840_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_839_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_838_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_837_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_836_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_835_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_834_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_833_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_832_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_831_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_830_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_829_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_828_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_827_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_826_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_825_sv2v_reg  <= w_data_i[0];
    end 
    if(N262) begin
      \xnz.mem_r_824_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_823_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_822_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_821_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_820_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_819_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_818_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_817_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_816_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_815_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_814_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_813_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_812_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_811_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_810_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_809_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_808_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_807_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_806_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_805_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_804_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_803_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_802_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_801_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_800_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_799_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_798_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_797_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_796_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_795_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_794_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_793_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_792_sv2v_reg  <= w_data_i[0];
    end 
    if(N261) begin
      \xnz.mem_r_791_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_790_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_789_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_788_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_787_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_786_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_785_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_784_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_783_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_782_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_781_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_780_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_779_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_778_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_777_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_776_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_775_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_774_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_773_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_772_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_771_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_770_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_769_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_768_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_767_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_766_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_765_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_764_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_763_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_762_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_761_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_760_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_759_sv2v_reg  <= w_data_i[0];
    end 
    if(N260) begin
      \xnz.mem_r_758_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_757_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_756_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_755_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_754_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_753_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_752_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_751_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_750_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_749_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_748_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_747_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_746_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_745_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_744_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_743_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_742_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_741_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_740_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_739_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_738_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_737_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_736_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_735_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_734_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_733_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_732_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_731_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_730_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_729_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_728_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_727_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_726_sv2v_reg  <= w_data_i[0];
    end 
    if(N259) begin
      \xnz.mem_r_725_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_724_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_723_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_722_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_721_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_720_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_719_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_718_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_717_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_716_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_715_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_714_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_713_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_712_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_711_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_710_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_709_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_708_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_707_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_706_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_705_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_704_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_703_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_702_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_701_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_700_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_699_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_698_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_697_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_696_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_695_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_694_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_693_sv2v_reg  <= w_data_i[0];
    end 
    if(N258) begin
      \xnz.mem_r_692_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_691_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_690_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_689_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_688_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_687_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_686_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_685_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_684_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_683_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_682_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_681_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_680_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_679_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_678_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_677_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_676_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_675_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_674_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_673_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_672_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_671_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_670_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_669_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_668_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_667_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_666_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_665_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_664_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_663_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_662_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_661_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_660_sv2v_reg  <= w_data_i[0];
    end 
    if(N257) begin
      \xnz.mem_r_659_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_658_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_657_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_656_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_655_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_654_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_653_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_652_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_651_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_650_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_649_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_648_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_647_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_646_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_645_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_644_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_643_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_642_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_641_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_640_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_639_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_638_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_637_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_636_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_635_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_634_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_633_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_632_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_631_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_630_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_629_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_628_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_627_sv2v_reg  <= w_data_i[0];
    end 
    if(N256) begin
      \xnz.mem_r_626_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_625_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_624_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_623_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_622_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_621_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_620_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_619_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_618_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_617_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_616_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_615_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_614_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_613_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_612_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_611_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_610_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_609_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_608_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_607_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_606_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_605_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_604_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_603_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_602_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_601_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_600_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_599_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_598_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_597_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_596_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_595_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_594_sv2v_reg  <= w_data_i[0];
    end 
    if(N255) begin
      \xnz.mem_r_593_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_592_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_591_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_590_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_589_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_588_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_587_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_586_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_585_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_584_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_583_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_582_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_581_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_580_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_579_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_578_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_577_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_576_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_575_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_574_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_573_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_572_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_571_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_570_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_569_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_568_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_567_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_566_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_565_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_564_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_563_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_562_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_561_sv2v_reg  <= w_data_i[0];
    end 
    if(N254) begin
      \xnz.mem_r_560_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_559_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_558_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_557_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_556_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_555_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_554_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_553_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_552_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_551_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_550_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_549_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_548_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_547_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_546_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_545_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_544_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_543_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_542_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_541_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_540_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_539_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_538_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_537_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_536_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_535_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_534_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_533_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_532_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_531_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_530_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_529_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_528_sv2v_reg  <= w_data_i[0];
    end 
    if(N253) begin
      \xnz.mem_r_527_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_526_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_525_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_524_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_523_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_522_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_521_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_520_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_519_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_518_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_517_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_516_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_515_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_514_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_513_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_512_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_511_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_510_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_509_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_508_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_507_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_506_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_505_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_504_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_503_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_502_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_501_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_500_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_499_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_498_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_497_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_496_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_495_sv2v_reg  <= w_data_i[0];
    end 
    if(N252) begin
      \xnz.mem_r_494_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_493_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_492_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_491_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_490_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_489_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_488_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_487_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_486_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_485_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_484_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_483_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_482_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_481_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_480_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_479_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_478_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_477_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_476_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_475_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_474_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_473_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_472_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_471_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_470_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_469_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_468_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_467_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_466_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_465_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_464_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_463_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_462_sv2v_reg  <= w_data_i[0];
    end 
    if(N251) begin
      \xnz.mem_r_461_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_460_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_459_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_458_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_457_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_456_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_455_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_454_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_453_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_452_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_451_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_450_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_449_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_448_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_447_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_446_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_445_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_444_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_443_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_442_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_441_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_440_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_439_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_438_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_437_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_436_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_435_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_434_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_433_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_432_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_431_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_430_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_429_sv2v_reg  <= w_data_i[0];
    end 
    if(N250) begin
      \xnz.mem_r_428_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_427_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_426_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_425_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_424_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_423_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_422_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_421_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_420_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_419_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_418_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_417_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_416_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_415_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_414_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_413_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_412_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_411_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_410_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_409_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_408_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_407_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_406_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_405_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_404_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_403_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_402_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_401_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_400_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_399_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_398_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_397_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_396_sv2v_reg  <= w_data_i[0];
    end 
    if(N249) begin
      \xnz.mem_r_395_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_394_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_393_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_392_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_391_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_390_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_389_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_388_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_387_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_386_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_385_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_384_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_383_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_382_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_381_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_380_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_379_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_378_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_377_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_376_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_375_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_374_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_373_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_372_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_371_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_370_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_369_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_368_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_367_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_366_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_365_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_364_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_363_sv2v_reg  <= w_data_i[0];
    end 
    if(N248) begin
      \xnz.mem_r_362_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_361_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_360_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_359_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_358_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_357_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_356_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_355_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_354_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_353_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_352_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_351_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_350_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_349_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_348_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_347_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_346_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_345_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_344_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_343_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_342_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_341_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_340_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_339_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_338_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_337_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_336_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_335_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_334_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_333_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_332_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_331_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_330_sv2v_reg  <= w_data_i[0];
    end 
    if(N247) begin
      \xnz.mem_r_329_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_328_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_327_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_326_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_325_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_324_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_323_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_322_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_321_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_320_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_319_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_318_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_317_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_316_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_315_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_314_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_313_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_312_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_311_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_310_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_309_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_308_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_307_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_306_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_305_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_304_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_303_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_302_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_301_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_300_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_299_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_298_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_297_sv2v_reg  <= w_data_i[0];
    end 
    if(N246) begin
      \xnz.mem_r_296_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_295_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_294_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_293_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_292_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_291_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_290_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_289_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_288_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_287_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_286_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_285_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_284_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_283_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_282_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_281_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_280_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_279_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_278_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_277_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_276_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_275_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_274_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_273_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_272_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_271_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_270_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_269_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_268_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_267_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_266_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_265_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_264_sv2v_reg  <= w_data_i[0];
    end 
    if(N245) begin
      \xnz.mem_r_263_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_262_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_261_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_260_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_259_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_258_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_257_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_256_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_255_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_254_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_253_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_252_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_251_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_250_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_249_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_248_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_247_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_246_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_245_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_244_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_243_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_242_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_241_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_240_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_239_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_238_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_237_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_236_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_235_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_234_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_233_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_232_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_231_sv2v_reg  <= w_data_i[0];
    end 
    if(N244) begin
      \xnz.mem_r_230_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_229_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_228_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_227_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_226_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_225_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_224_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_223_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_222_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_221_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_220_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_219_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_218_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_217_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_216_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_215_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_214_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_213_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_212_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_211_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_210_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_209_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_208_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_207_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_206_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_205_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_204_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_203_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_202_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_201_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_200_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_199_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_198_sv2v_reg  <= w_data_i[0];
    end 
    if(N243) begin
      \xnz.mem_r_197_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_196_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_195_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_194_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_193_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_192_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_191_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_190_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_189_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_188_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_187_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_186_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_185_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_184_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_183_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_182_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_181_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_180_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_179_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_178_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_177_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_176_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_175_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_174_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_173_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_172_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_171_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_170_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_169_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_168_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_167_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_166_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_165_sv2v_reg  <= w_data_i[0];
    end 
    if(N242) begin
      \xnz.mem_r_164_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_163_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_162_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_161_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_160_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_159_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_158_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_157_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_156_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_155_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_154_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_153_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_152_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_151_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_150_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_149_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_148_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_147_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_146_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_145_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_144_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_143_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_142_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_141_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_140_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_139_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_138_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_137_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_136_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_135_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_134_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_133_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_132_sv2v_reg  <= w_data_i[0];
    end 
    if(N241) begin
      \xnz.mem_r_131_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_130_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_129_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_128_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_127_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_126_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_125_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_124_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_123_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_122_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_121_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_120_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_119_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_118_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_117_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_116_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_115_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_114_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_113_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_112_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_111_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_110_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_109_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_108_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_107_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_106_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_105_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_104_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_103_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_102_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_101_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_100_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_99_sv2v_reg  <= w_data_i[0];
    end 
    if(N240) begin
      \xnz.mem_r_98_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_97_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_96_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_95_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_94_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_93_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_92_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_91_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_90_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_89_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_88_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_87_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_86_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_85_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_84_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_83_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_82_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_81_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_80_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_79_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_78_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_77_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_76_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_75_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_74_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_73_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_72_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_71_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_70_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_69_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_68_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_67_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_66_sv2v_reg  <= w_data_i[0];
    end 
    if(N239) begin
      \xnz.mem_r_65_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_64_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_63_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_62_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_61_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_60_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_59_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_58_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_57_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_56_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_55_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_54_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_53_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_52_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_51_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_50_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_49_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_48_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_47_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_46_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_45_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_44_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_43_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_42_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_41_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_40_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_39_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_38_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_37_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_36_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_35_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_34_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_33_sv2v_reg  <= w_data_i[0];
    end 
    if(N238) begin
      \xnz.mem_r_32_sv2v_reg  <= w_data_i[32];
      \xnz.mem_r_31_sv2v_reg  <= w_data_i[31];
      \xnz.mem_r_30_sv2v_reg  <= w_data_i[30];
      \xnz.mem_r_29_sv2v_reg  <= w_data_i[29];
      \xnz.mem_r_28_sv2v_reg  <= w_data_i[28];
      \xnz.mem_r_27_sv2v_reg  <= w_data_i[27];
      \xnz.mem_r_26_sv2v_reg  <= w_data_i[26];
      \xnz.mem_r_25_sv2v_reg  <= w_data_i[25];
      \xnz.mem_r_24_sv2v_reg  <= w_data_i[24];
      \xnz.mem_r_23_sv2v_reg  <= w_data_i[23];
      \xnz.mem_r_22_sv2v_reg  <= w_data_i[22];
      \xnz.mem_r_21_sv2v_reg  <= w_data_i[21];
      \xnz.mem_r_20_sv2v_reg  <= w_data_i[20];
      \xnz.mem_r_19_sv2v_reg  <= w_data_i[19];
      \xnz.mem_r_18_sv2v_reg  <= w_data_i[18];
      \xnz.mem_r_17_sv2v_reg  <= w_data_i[17];
      \xnz.mem_r_16_sv2v_reg  <= w_data_i[16];
      \xnz.mem_r_15_sv2v_reg  <= w_data_i[15];
      \xnz.mem_r_14_sv2v_reg  <= w_data_i[14];
      \xnz.mem_r_13_sv2v_reg  <= w_data_i[13];
      \xnz.mem_r_12_sv2v_reg  <= w_data_i[12];
      \xnz.mem_r_11_sv2v_reg  <= w_data_i[11];
      \xnz.mem_r_10_sv2v_reg  <= w_data_i[10];
      \xnz.mem_r_9_sv2v_reg  <= w_data_i[9];
      \xnz.mem_r_8_sv2v_reg  <= w_data_i[8];
      \xnz.mem_r_7_sv2v_reg  <= w_data_i[7];
      \xnz.mem_r_6_sv2v_reg  <= w_data_i[6];
      \xnz.mem_r_5_sv2v_reg  <= w_data_i[5];
      \xnz.mem_r_4_sv2v_reg  <= w_data_i[4];
      \xnz.mem_r_3_sv2v_reg  <= w_data_i[3];
      \xnz.mem_r_2_sv2v_reg  <= w_data_i[2];
      \xnz.mem_r_1_sv2v_reg  <= w_data_i[1];
      \xnz.mem_r_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module regfile_width_p33_els_p32_num_rs_p3_x0_tied_to_zero_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [4:0] w_addr_i;
  input [32:0] w_data_i;
  input [2:0] r_v_i;
  input [14:0] r_addr_i;
  output [98:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  wire [98:0] r_data_o;

  regfile_synth_width_p33_els_p32_num_rs_p3_x0_tied_to_zero_p0
  \synth.rf 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_transpose_width_p3_els_p1
(
  i,
  o
);

  input [2:0] i;
  output [2:0] o;
  wire [2:0] o;
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module scoreboard_els_p32_num_src_port_p3_num_clear_port_p1_x0_tied_to_zero_p0
(
  clk_i,
  reset_i,
  src_id_i,
  dest_id_i,
  op_reads_rf_i,
  op_writes_rf_i,
  score_i,
  score_id_i,
  clear_i,
  clear_id_i,
  dependency_o
);

  input [14:0] src_id_i;
  input [4:0] dest_id_i;
  input [2:0] op_reads_rf_i;
  input [4:0] score_id_i;
  input [0:0] clear_i;
  input [4:0] clear_id_i;
  input clk_i;
  input reset_i;
  input op_writes_rf_i;
  input score_i;
  output dependency_o;
  wire dependency_o,_0_net_,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,rd_depend_on_sb,N264,N265,N266,N267,N268,N269,
  N270,N271,rd_depend_on_score,depend_on_sb,depend_on_score,N272,N273,N274,N275,N276,
  N277,N278,N279,N280,N281,N282,N283,N284,N285;
  wire [31:0] clear_by_port,clear_by_port_t,score_bits,scoreboard_r;
  wire [2:0] rs_depend_on_sb,rs_on_clear,rs_on_clear_t,rs_depend_on_score;
  wire [0:0] rd_on_clear;
  reg scoreboard_r_31_sv2v_reg,scoreboard_r_30_sv2v_reg,scoreboard_r_29_sv2v_reg,
  scoreboard_r_28_sv2v_reg,scoreboard_r_27_sv2v_reg,scoreboard_r_26_sv2v_reg,
  scoreboard_r_25_sv2v_reg,scoreboard_r_24_sv2v_reg,scoreboard_r_23_sv2v_reg,
  scoreboard_r_22_sv2v_reg,scoreboard_r_21_sv2v_reg,scoreboard_r_20_sv2v_reg,
  scoreboard_r_19_sv2v_reg,scoreboard_r_18_sv2v_reg,scoreboard_r_17_sv2v_reg,scoreboard_r_16_sv2v_reg,
  scoreboard_r_15_sv2v_reg,scoreboard_r_14_sv2v_reg,scoreboard_r_13_sv2v_reg,
  scoreboard_r_12_sv2v_reg,scoreboard_r_11_sv2v_reg,scoreboard_r_10_sv2v_reg,
  scoreboard_r_9_sv2v_reg,scoreboard_r_8_sv2v_reg,scoreboard_r_7_sv2v_reg,
  scoreboard_r_6_sv2v_reg,scoreboard_r_5_sv2v_reg,scoreboard_r_4_sv2v_reg,scoreboard_r_3_sv2v_reg,
  scoreboard_r_2_sv2v_reg,scoreboard_r_1_sv2v_reg,scoreboard_r_0_sv2v_reg;
  assign scoreboard_r[31] = scoreboard_r_31_sv2v_reg;
  assign scoreboard_r[30] = scoreboard_r_30_sv2v_reg;
  assign scoreboard_r[29] = scoreboard_r_29_sv2v_reg;
  assign scoreboard_r[28] = scoreboard_r_28_sv2v_reg;
  assign scoreboard_r[27] = scoreboard_r_27_sv2v_reg;
  assign scoreboard_r[26] = scoreboard_r_26_sv2v_reg;
  assign scoreboard_r[25] = scoreboard_r_25_sv2v_reg;
  assign scoreboard_r[24] = scoreboard_r_24_sv2v_reg;
  assign scoreboard_r[23] = scoreboard_r_23_sv2v_reg;
  assign scoreboard_r[22] = scoreboard_r_22_sv2v_reg;
  assign scoreboard_r[21] = scoreboard_r_21_sv2v_reg;
  assign scoreboard_r[20] = scoreboard_r_20_sv2v_reg;
  assign scoreboard_r[19] = scoreboard_r_19_sv2v_reg;
  assign scoreboard_r[18] = scoreboard_r_18_sv2v_reg;
  assign scoreboard_r[17] = scoreboard_r_17_sv2v_reg;
  assign scoreboard_r[16] = scoreboard_r_16_sv2v_reg;
  assign scoreboard_r[15] = scoreboard_r_15_sv2v_reg;
  assign scoreboard_r[14] = scoreboard_r_14_sv2v_reg;
  assign scoreboard_r[13] = scoreboard_r_13_sv2v_reg;
  assign scoreboard_r[12] = scoreboard_r_12_sv2v_reg;
  assign scoreboard_r[11] = scoreboard_r_11_sv2v_reg;
  assign scoreboard_r[10] = scoreboard_r_10_sv2v_reg;
  assign scoreboard_r[9] = scoreboard_r_9_sv2v_reg;
  assign scoreboard_r[8] = scoreboard_r_8_sv2v_reg;
  assign scoreboard_r[7] = scoreboard_r_7_sv2v_reg;
  assign scoreboard_r[6] = scoreboard_r_6_sv2v_reg;
  assign scoreboard_r[5] = scoreboard_r_5_sv2v_reg;
  assign scoreboard_r[4] = scoreboard_r_4_sv2v_reg;
  assign scoreboard_r[3] = scoreboard_r_3_sv2v_reg;
  assign scoreboard_r[2] = scoreboard_r_2_sv2v_reg;
  assign scoreboard_r[1] = scoreboard_r_1_sv2v_reg;
  assign scoreboard_r[0] = scoreboard_r_0_sv2v_reg;

  bsg_transpose_width_p32_els_p1
  tranposer
  (
    .i(clear_by_port),
    .o(clear_by_port_t)
  );


  bsg_decode_with_v_num_out_p32
  \clr_dcode_v_0_.clear_decode_v 
  (
    .i(clear_id_i),
    .v_i(clear_i[0]),
    .o(clear_by_port)
  );


  bsg_decode_with_v_num_out_p32
  score_demux
  (
    .i(score_id_i),
    .v_i(_0_net_),
    .o(score_bits)
  );

  assign N65 = (N33)? scoreboard_r[0] : 
               (N35)? scoreboard_r[1] : 
               (N37)? scoreboard_r[2] : 
               (N39)? scoreboard_r[3] : 
               (N41)? scoreboard_r[4] : 
               (N43)? scoreboard_r[5] : 
               (N45)? scoreboard_r[6] : 
               (N47)? scoreboard_r[7] : 
               (N49)? scoreboard_r[8] : 
               (N51)? scoreboard_r[9] : 
               (N53)? scoreboard_r[10] : 
               (N55)? scoreboard_r[11] : 
               (N57)? scoreboard_r[12] : 
               (N59)? scoreboard_r[13] : 
               (N61)? scoreboard_r[14] : 
               (N63)? scoreboard_r[15] : 
               (N34)? scoreboard_r[16] : 
               (N36)? scoreboard_r[17] : 
               (N38)? scoreboard_r[18] : 
               (N40)? scoreboard_r[19] : 
               (N42)? scoreboard_r[20] : 
               (N44)? scoreboard_r[21] : 
               (N46)? scoreboard_r[22] : 
               (N48)? scoreboard_r[23] : 
               (N50)? scoreboard_r[24] : 
               (N52)? scoreboard_r[25] : 
               (N54)? scoreboard_r[26] : 
               (N56)? scoreboard_r[27] : 
               (N58)? scoreboard_r[28] : 
               (N60)? scoreboard_r[29] : 
               (N62)? scoreboard_r[30] : 
               (N64)? scoreboard_r[31] : 1'b0;
  assign N131 = (N99)? scoreboard_r[0] : 
                (N101)? scoreboard_r[1] : 
                (N103)? scoreboard_r[2] : 
                (N105)? scoreboard_r[3] : 
                (N107)? scoreboard_r[4] : 
                (N109)? scoreboard_r[5] : 
                (N111)? scoreboard_r[6] : 
                (N113)? scoreboard_r[7] : 
                (N115)? scoreboard_r[8] : 
                (N117)? scoreboard_r[9] : 
                (N119)? scoreboard_r[10] : 
                (N121)? scoreboard_r[11] : 
                (N123)? scoreboard_r[12] : 
                (N125)? scoreboard_r[13] : 
                (N127)? scoreboard_r[14] : 
                (N129)? scoreboard_r[15] : 
                (N100)? scoreboard_r[16] : 
                (N102)? scoreboard_r[17] : 
                (N104)? scoreboard_r[18] : 
                (N106)? scoreboard_r[19] : 
                (N108)? scoreboard_r[20] : 
                (N110)? scoreboard_r[21] : 
                (N112)? scoreboard_r[22] : 
                (N114)? scoreboard_r[23] : 
                (N116)? scoreboard_r[24] : 
                (N118)? scoreboard_r[25] : 
                (N120)? scoreboard_r[26] : 
                (N122)? scoreboard_r[27] : 
                (N124)? scoreboard_r[28] : 
                (N126)? scoreboard_r[29] : 
                (N128)? scoreboard_r[30] : 
                (N130)? scoreboard_r[31] : 1'b0;
  assign N197 = (N165)? scoreboard_r[0] : 
                (N167)? scoreboard_r[1] : 
                (N169)? scoreboard_r[2] : 
                (N171)? scoreboard_r[3] : 
                (N173)? scoreboard_r[4] : 
                (N175)? scoreboard_r[5] : 
                (N177)? scoreboard_r[6] : 
                (N179)? scoreboard_r[7] : 
                (N181)? scoreboard_r[8] : 
                (N183)? scoreboard_r[9] : 
                (N185)? scoreboard_r[10] : 
                (N187)? scoreboard_r[11] : 
                (N189)? scoreboard_r[12] : 
                (N191)? scoreboard_r[13] : 
                (N193)? scoreboard_r[14] : 
                (N195)? scoreboard_r[15] : 
                (N166)? scoreboard_r[16] : 
                (N168)? scoreboard_r[17] : 
                (N170)? scoreboard_r[18] : 
                (N172)? scoreboard_r[19] : 
                (N174)? scoreboard_r[20] : 
                (N176)? scoreboard_r[21] : 
                (N178)? scoreboard_r[22] : 
                (N180)? scoreboard_r[23] : 
                (N182)? scoreboard_r[24] : 
                (N184)? scoreboard_r[25] : 
                (N186)? scoreboard_r[26] : 
                (N188)? scoreboard_r[27] : 
                (N190)? scoreboard_r[28] : 
                (N192)? scoreboard_r[29] : 
                (N194)? scoreboard_r[30] : 
                (N196)? scoreboard_r[31] : 1'b0;
  assign N263 = (N231)? scoreboard_r[0] : 
                (N233)? scoreboard_r[1] : 
                (N235)? scoreboard_r[2] : 
                (N237)? scoreboard_r[3] : 
                (N239)? scoreboard_r[4] : 
                (N241)? scoreboard_r[5] : 
                (N243)? scoreboard_r[6] : 
                (N245)? scoreboard_r[7] : 
                (N247)? scoreboard_r[8] : 
                (N249)? scoreboard_r[9] : 
                (N251)? scoreboard_r[10] : 
                (N253)? scoreboard_r[11] : 
                (N255)? scoreboard_r[12] : 
                (N257)? scoreboard_r[13] : 
                (N259)? scoreboard_r[14] : 
                (N261)? scoreboard_r[15] : 
                (N232)? scoreboard_r[16] : 
                (N234)? scoreboard_r[17] : 
                (N236)? scoreboard_r[18] : 
                (N238)? scoreboard_r[19] : 
                (N240)? scoreboard_r[20] : 
                (N242)? scoreboard_r[21] : 
                (N244)? scoreboard_r[22] : 
                (N246)? scoreboard_r[23] : 
                (N248)? scoreboard_r[24] : 
                (N250)? scoreboard_r[25] : 
                (N252)? scoreboard_r[26] : 
                (N254)? scoreboard_r[27] : 
                (N256)? scoreboard_r[28] : 
                (N258)? scoreboard_r[29] : 
                (N260)? scoreboard_r[30] : 
                (N262)? scoreboard_r[31] : 1'b0;
  assign N264 = clear_id_i == src_id_i[4:0];
  assign N265 = clear_id_i == src_id_i[9:5];
  assign N266 = clear_id_i == src_id_i[14:10];
  assign N267 = clear_id_i == dest_id_i;

  bsg_transpose_width_p3_els_p1
  trans1
  (
    .i(rs_on_clear),
    .o(rs_on_clear_t)
  );

  assign N268 = src_id_i[4:0] == score_id_i;
  assign N269 = src_id_i[9:5] == score_id_i;
  assign N270 = src_id_i[14:10] == score_id_i;
  assign N271 = dest_id_i == score_id_i;
  assign _0_net_ = score_i & 1'b1;
  assign N0 = ~src_id_i[0];
  assign N1 = ~src_id_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & src_id_i[1];
  assign N4 = src_id_i[0] & N1;
  assign N5 = src_id_i[0] & src_id_i[1];
  assign N6 = ~src_id_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & src_id_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & src_id_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & src_id_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & src_id_i[2];
  assign N15 = ~src_id_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & src_id_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & src_id_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & src_id_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & src_id_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & src_id_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & src_id_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & src_id_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & src_id_i[3];
  assign N32 = ~src_id_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & src_id_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & src_id_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & src_id_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & src_id_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & src_id_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & src_id_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & src_id_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & src_id_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & src_id_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & src_id_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & src_id_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & src_id_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & src_id_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & src_id_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & src_id_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & src_id_i[4];
  assign rs_depend_on_sb[0] = N65 & op_reads_rf_i[0];
  assign N66 = ~src_id_i[5];
  assign N67 = ~src_id_i[6];
  assign N68 = N66 & N67;
  assign N69 = N66 & src_id_i[6];
  assign N70 = src_id_i[5] & N67;
  assign N71 = src_id_i[5] & src_id_i[6];
  assign N72 = ~src_id_i[7];
  assign N73 = N68 & N72;
  assign N74 = N68 & src_id_i[7];
  assign N75 = N70 & N72;
  assign N76 = N70 & src_id_i[7];
  assign N77 = N69 & N72;
  assign N78 = N69 & src_id_i[7];
  assign N79 = N71 & N72;
  assign N80 = N71 & src_id_i[7];
  assign N81 = ~src_id_i[8];
  assign N82 = N73 & N81;
  assign N83 = N73 & src_id_i[8];
  assign N84 = N75 & N81;
  assign N85 = N75 & src_id_i[8];
  assign N86 = N77 & N81;
  assign N87 = N77 & src_id_i[8];
  assign N88 = N79 & N81;
  assign N89 = N79 & src_id_i[8];
  assign N90 = N74 & N81;
  assign N91 = N74 & src_id_i[8];
  assign N92 = N76 & N81;
  assign N93 = N76 & src_id_i[8];
  assign N94 = N78 & N81;
  assign N95 = N78 & src_id_i[8];
  assign N96 = N80 & N81;
  assign N97 = N80 & src_id_i[8];
  assign N98 = ~src_id_i[9];
  assign N99 = N82 & N98;
  assign N100 = N82 & src_id_i[9];
  assign N101 = N84 & N98;
  assign N102 = N84 & src_id_i[9];
  assign N103 = N86 & N98;
  assign N104 = N86 & src_id_i[9];
  assign N105 = N88 & N98;
  assign N106 = N88 & src_id_i[9];
  assign N107 = N90 & N98;
  assign N108 = N90 & src_id_i[9];
  assign N109 = N92 & N98;
  assign N110 = N92 & src_id_i[9];
  assign N111 = N94 & N98;
  assign N112 = N94 & src_id_i[9];
  assign N113 = N96 & N98;
  assign N114 = N96 & src_id_i[9];
  assign N115 = N83 & N98;
  assign N116 = N83 & src_id_i[9];
  assign N117 = N85 & N98;
  assign N118 = N85 & src_id_i[9];
  assign N119 = N87 & N98;
  assign N120 = N87 & src_id_i[9];
  assign N121 = N89 & N98;
  assign N122 = N89 & src_id_i[9];
  assign N123 = N91 & N98;
  assign N124 = N91 & src_id_i[9];
  assign N125 = N93 & N98;
  assign N126 = N93 & src_id_i[9];
  assign N127 = N95 & N98;
  assign N128 = N95 & src_id_i[9];
  assign N129 = N97 & N98;
  assign N130 = N97 & src_id_i[9];
  assign rs_depend_on_sb[1] = N131 & op_reads_rf_i[1];
  assign N132 = ~src_id_i[10];
  assign N133 = ~src_id_i[11];
  assign N134 = N132 & N133;
  assign N135 = N132 & src_id_i[11];
  assign N136 = src_id_i[10] & N133;
  assign N137 = src_id_i[10] & src_id_i[11];
  assign N138 = ~src_id_i[12];
  assign N139 = N134 & N138;
  assign N140 = N134 & src_id_i[12];
  assign N141 = N136 & N138;
  assign N142 = N136 & src_id_i[12];
  assign N143 = N135 & N138;
  assign N144 = N135 & src_id_i[12];
  assign N145 = N137 & N138;
  assign N146 = N137 & src_id_i[12];
  assign N147 = ~src_id_i[13];
  assign N148 = N139 & N147;
  assign N149 = N139 & src_id_i[13];
  assign N150 = N141 & N147;
  assign N151 = N141 & src_id_i[13];
  assign N152 = N143 & N147;
  assign N153 = N143 & src_id_i[13];
  assign N154 = N145 & N147;
  assign N155 = N145 & src_id_i[13];
  assign N156 = N140 & N147;
  assign N157 = N140 & src_id_i[13];
  assign N158 = N142 & N147;
  assign N159 = N142 & src_id_i[13];
  assign N160 = N144 & N147;
  assign N161 = N144 & src_id_i[13];
  assign N162 = N146 & N147;
  assign N163 = N146 & src_id_i[13];
  assign N164 = ~src_id_i[14];
  assign N165 = N148 & N164;
  assign N166 = N148 & src_id_i[14];
  assign N167 = N150 & N164;
  assign N168 = N150 & src_id_i[14];
  assign N169 = N152 & N164;
  assign N170 = N152 & src_id_i[14];
  assign N171 = N154 & N164;
  assign N172 = N154 & src_id_i[14];
  assign N173 = N156 & N164;
  assign N174 = N156 & src_id_i[14];
  assign N175 = N158 & N164;
  assign N176 = N158 & src_id_i[14];
  assign N177 = N160 & N164;
  assign N178 = N160 & src_id_i[14];
  assign N179 = N162 & N164;
  assign N180 = N162 & src_id_i[14];
  assign N181 = N149 & N164;
  assign N182 = N149 & src_id_i[14];
  assign N183 = N151 & N164;
  assign N184 = N151 & src_id_i[14];
  assign N185 = N153 & N164;
  assign N186 = N153 & src_id_i[14];
  assign N187 = N155 & N164;
  assign N188 = N155 & src_id_i[14];
  assign N189 = N157 & N164;
  assign N190 = N157 & src_id_i[14];
  assign N191 = N159 & N164;
  assign N192 = N159 & src_id_i[14];
  assign N193 = N161 & N164;
  assign N194 = N161 & src_id_i[14];
  assign N195 = N163 & N164;
  assign N196 = N163 & src_id_i[14];
  assign rs_depend_on_sb[2] = N197 & op_reads_rf_i[2];
  assign N198 = ~dest_id_i[0];
  assign N199 = ~dest_id_i[1];
  assign N200 = N198 & N199;
  assign N201 = N198 & dest_id_i[1];
  assign N202 = dest_id_i[0] & N199;
  assign N203 = dest_id_i[0] & dest_id_i[1];
  assign N204 = ~dest_id_i[2];
  assign N205 = N200 & N204;
  assign N206 = N200 & dest_id_i[2];
  assign N207 = N202 & N204;
  assign N208 = N202 & dest_id_i[2];
  assign N209 = N201 & N204;
  assign N210 = N201 & dest_id_i[2];
  assign N211 = N203 & N204;
  assign N212 = N203 & dest_id_i[2];
  assign N213 = ~dest_id_i[3];
  assign N214 = N205 & N213;
  assign N215 = N205 & dest_id_i[3];
  assign N216 = N207 & N213;
  assign N217 = N207 & dest_id_i[3];
  assign N218 = N209 & N213;
  assign N219 = N209 & dest_id_i[3];
  assign N220 = N211 & N213;
  assign N221 = N211 & dest_id_i[3];
  assign N222 = N206 & N213;
  assign N223 = N206 & dest_id_i[3];
  assign N224 = N208 & N213;
  assign N225 = N208 & dest_id_i[3];
  assign N226 = N210 & N213;
  assign N227 = N210 & dest_id_i[3];
  assign N228 = N212 & N213;
  assign N229 = N212 & dest_id_i[3];
  assign N230 = ~dest_id_i[4];
  assign N231 = N214 & N230;
  assign N232 = N214 & dest_id_i[4];
  assign N233 = N216 & N230;
  assign N234 = N216 & dest_id_i[4];
  assign N235 = N218 & N230;
  assign N236 = N218 & dest_id_i[4];
  assign N237 = N220 & N230;
  assign N238 = N220 & dest_id_i[4];
  assign N239 = N222 & N230;
  assign N240 = N222 & dest_id_i[4];
  assign N241 = N224 & N230;
  assign N242 = N224 & dest_id_i[4];
  assign N243 = N226 & N230;
  assign N244 = N226 & dest_id_i[4];
  assign N245 = N228 & N230;
  assign N246 = N228 & dest_id_i[4];
  assign N247 = N215 & N230;
  assign N248 = N215 & dest_id_i[4];
  assign N249 = N217 & N230;
  assign N250 = N217 & dest_id_i[4];
  assign N251 = N219 & N230;
  assign N252 = N219 & dest_id_i[4];
  assign N253 = N221 & N230;
  assign N254 = N221 & dest_id_i[4];
  assign N255 = N223 & N230;
  assign N256 = N223 & dest_id_i[4];
  assign N257 = N225 & N230;
  assign N258 = N225 & dest_id_i[4];
  assign N259 = N227 & N230;
  assign N260 = N227 & dest_id_i[4];
  assign N261 = N229 & N230;
  assign N262 = N229 & dest_id_i[4];
  assign rd_depend_on_sb = N263 & op_writes_rf_i;
  assign rs_on_clear[0] = clear_i[0] & N264;
  assign rs_on_clear[1] = clear_i[0] & N265;
  assign rs_on_clear[2] = clear_i[0] & N266;
  assign rd_on_clear[0] = clear_i[0] & N267;
  assign rs_depend_on_score[0] = N268 & op_reads_rf_i[0];
  assign rs_depend_on_score[1] = N269 & op_reads_rf_i[1];
  assign rs_depend_on_score[2] = N270 & op_reads_rf_i[2];
  assign rd_depend_on_score = N271 & op_writes_rf_i;
  assign depend_on_sb = N279 | N281;
  assign N279 = N276 | N278;
  assign N276 = N273 | N275;
  assign N273 = rd_depend_on_sb & N272;
  assign N272 = ~rd_on_clear[0];
  assign N275 = rs_depend_on_sb[2] & N274;
  assign N274 = ~rs_on_clear_t[2];
  assign N278 = rs_depend_on_sb[1] & N277;
  assign N277 = ~rs_on_clear_t[1];
  assign N281 = rs_depend_on_sb[0] & N280;
  assign N280 = ~rs_on_clear_t[0];
  assign depend_on_score = N283 | rs_depend_on_score[0];
  assign N283 = N282 | rs_depend_on_score[1];
  assign N282 = rd_depend_on_score | rs_depend_on_score[2];
  assign dependency_o = depend_on_sb | N285;
  assign N285 = N284 & 1'b1;
  assign N284 = depend_on_score & score_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      scoreboard_r_31_sv2v_reg <= 1'b0;
    end else if(score_bits[31]) begin
      scoreboard_r_31_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[31]) begin
      scoreboard_r_31_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_30_sv2v_reg <= 1'b0;
    end else if(score_bits[30]) begin
      scoreboard_r_30_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[30]) begin
      scoreboard_r_30_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_29_sv2v_reg <= 1'b0;
    end else if(score_bits[29]) begin
      scoreboard_r_29_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[29]) begin
      scoreboard_r_29_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_28_sv2v_reg <= 1'b0;
    end else if(score_bits[28]) begin
      scoreboard_r_28_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[28]) begin
      scoreboard_r_28_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_27_sv2v_reg <= 1'b0;
    end else if(score_bits[27]) begin
      scoreboard_r_27_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[27]) begin
      scoreboard_r_27_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_26_sv2v_reg <= 1'b0;
    end else if(score_bits[26]) begin
      scoreboard_r_26_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[26]) begin
      scoreboard_r_26_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_25_sv2v_reg <= 1'b0;
    end else if(score_bits[25]) begin
      scoreboard_r_25_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[25]) begin
      scoreboard_r_25_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_24_sv2v_reg <= 1'b0;
    end else if(score_bits[24]) begin
      scoreboard_r_24_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[24]) begin
      scoreboard_r_24_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_23_sv2v_reg <= 1'b0;
    end else if(score_bits[23]) begin
      scoreboard_r_23_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[23]) begin
      scoreboard_r_23_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_22_sv2v_reg <= 1'b0;
    end else if(score_bits[22]) begin
      scoreboard_r_22_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[22]) begin
      scoreboard_r_22_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_21_sv2v_reg <= 1'b0;
    end else if(score_bits[21]) begin
      scoreboard_r_21_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[21]) begin
      scoreboard_r_21_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_20_sv2v_reg <= 1'b0;
    end else if(score_bits[20]) begin
      scoreboard_r_20_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[20]) begin
      scoreboard_r_20_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_19_sv2v_reg <= 1'b0;
    end else if(score_bits[19]) begin
      scoreboard_r_19_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[19]) begin
      scoreboard_r_19_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_18_sv2v_reg <= 1'b0;
    end else if(score_bits[18]) begin
      scoreboard_r_18_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[18]) begin
      scoreboard_r_18_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_17_sv2v_reg <= 1'b0;
    end else if(score_bits[17]) begin
      scoreboard_r_17_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[17]) begin
      scoreboard_r_17_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_16_sv2v_reg <= 1'b0;
    end else if(score_bits[16]) begin
      scoreboard_r_16_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[16]) begin
      scoreboard_r_16_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_15_sv2v_reg <= 1'b0;
    end else if(score_bits[15]) begin
      scoreboard_r_15_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[15]) begin
      scoreboard_r_15_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_14_sv2v_reg <= 1'b0;
    end else if(score_bits[14]) begin
      scoreboard_r_14_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[14]) begin
      scoreboard_r_14_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_13_sv2v_reg <= 1'b0;
    end else if(score_bits[13]) begin
      scoreboard_r_13_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[13]) begin
      scoreboard_r_13_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_12_sv2v_reg <= 1'b0;
    end else if(score_bits[12]) begin
      scoreboard_r_12_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[12]) begin
      scoreboard_r_12_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_11_sv2v_reg <= 1'b0;
    end else if(score_bits[11]) begin
      scoreboard_r_11_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[11]) begin
      scoreboard_r_11_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_10_sv2v_reg <= 1'b0;
    end else if(score_bits[10]) begin
      scoreboard_r_10_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[10]) begin
      scoreboard_r_10_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_9_sv2v_reg <= 1'b0;
    end else if(score_bits[9]) begin
      scoreboard_r_9_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[9]) begin
      scoreboard_r_9_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_8_sv2v_reg <= 1'b0;
    end else if(score_bits[8]) begin
      scoreboard_r_8_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[8]) begin
      scoreboard_r_8_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_7_sv2v_reg <= 1'b0;
    end else if(score_bits[7]) begin
      scoreboard_r_7_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[7]) begin
      scoreboard_r_7_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_6_sv2v_reg <= 1'b0;
    end else if(score_bits[6]) begin
      scoreboard_r_6_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[6]) begin
      scoreboard_r_6_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_5_sv2v_reg <= 1'b0;
    end else if(score_bits[5]) begin
      scoreboard_r_5_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[5]) begin
      scoreboard_r_5_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_4_sv2v_reg <= 1'b0;
    end else if(score_bits[4]) begin
      scoreboard_r_4_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[4]) begin
      scoreboard_r_4_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_3_sv2v_reg <= 1'b0;
    end else if(score_bits[3]) begin
      scoreboard_r_3_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[3]) begin
      scoreboard_r_3_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_2_sv2v_reg <= 1'b0;
    end else if(score_bits[2]) begin
      scoreboard_r_2_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[2]) begin
      scoreboard_r_2_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_1_sv2v_reg <= 1'b0;
    end else if(score_bits[1]) begin
      scoreboard_r_1_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[1]) begin
      scoreboard_r_1_sv2v_reg <= 1'b0;
    end 
    if(reset_i) begin
      scoreboard_r_0_sv2v_reg <= 1'b0;
    end else if(score_bits[0]) begin
      scoreboard_r_0_sv2v_reg <= 1'b1;
    end else if(clear_by_port_t[0]) begin
      scoreboard_r_0_sv2v_reg <= 1'b0;
    end 
  end


endmodule



module fcsr
(
  clk_i,
  reset_i,
  v_i,
  funct3_i,
  rs1_i,
  data_i,
  addr_i,
  data_o,
  data_v_o,
  fflags_v_i,
  fflags_i,
  frm_o
);

  input [2:0] funct3_i;
  input [4:0] rs1_i;
  input [7:0] data_i;
  input [11:0] addr_i;
  output [7:0] data_o;
  input [1:0] fflags_v_i;
  input [9:0] fflags_i;
  output [2:0] frm_o;
  input clk_i;
  input reset_i;
  input v_i;
  output data_v_o;
  wire [7:0] data_o,write_mask,write_data;
  wire [2:0] frm_o,frm_write_mask,frm_write_data;
  wire data_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135;
  wire [9:0] filtered_fflags;
  wire [4:0] combined_fflags,fflags_write_mask,fflags_write_data,fflags_r;
  reg fflags_r_4_sv2v_reg,fflags_r_3_sv2v_reg,fflags_r_2_sv2v_reg,fflags_r_1_sv2v_reg,
  fflags_r_0_sv2v_reg,frm_o_2_sv2v_reg,frm_o_1_sv2v_reg,frm_o_0_sv2v_reg;
  assign fflags_r[4] = fflags_r_4_sv2v_reg;
  assign fflags_r[3] = fflags_r_3_sv2v_reg;
  assign fflags_r[2] = fflags_r_2_sv2v_reg;
  assign fflags_r[1] = fflags_r_1_sv2v_reg;
  assign fflags_r[0] = fflags_r_0_sv2v_reg;
  assign frm_o[2] = frm_o_2_sv2v_reg;
  assign frm_o[1] = frm_o_1_sv2v_reg;
  assign frm_o[0] = frm_o_0_sv2v_reg;
  assign N19 = funct3_i[2] | funct3_i[1];
  assign N20 = N19 | N37;
  assign N22 = funct3_i[2] | N36;
  assign N23 = N22 | funct3_i[0];
  assign N25 = N22 | N37;
  assign N28 = N27 | funct3_i[1];
  assign N29 = N28 | N37;
  assign N31 = N27 | N36;
  assign N32 = N31 | funct3_i[0];
  assign N34 = funct3_i[2] & funct3_i[1];
  assign N35 = N34 & funct3_i[0];
  assign N38 = N36 & N37;
  assign N68 = addr_i[11] | addr_i[10];
  assign N69 = addr_i[9] | addr_i[8];
  assign N70 = addr_i[7] | addr_i[6];
  assign N71 = addr_i[5] | addr_i[4];
  assign N72 = addr_i[3] | addr_i[2];
  assign N73 = N68 | N69;
  assign N74 = N70 | N71;
  assign N75 = N72 | N124;
  assign N76 = N73 | N74;
  assign N77 = N76 | N75;
  assign N86 = N113 & addr_i[0];
  assign N87 = N116 & N86;
  assign N109 = N99 & N100;
  assign N110 = N101 & N102;
  assign N111 = N103 & N104;
  assign N112 = N105 & N106;
  assign N113 = N107 & N108;
  assign N114 = N109 & N110;
  assign N115 = N111 & N112;
  assign N116 = N114 & N115;
  assign N117 = N116 & N113;
  assign N119 = addr_i[1] | N125;
  assign N121 = N124 | addr_i[0];
  assign N123 = addr_i[1] & addr_i[0];
  assign N126 = N124 & N125;
  assign { N59, N58, N57, N56, N55, N54, N53, N52 } = (N0)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                      (N1)? data_i : 
                                                      (N2)? data_i : 
                                                      (N3)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                      (N4)? { 1'b0, 1'b0, 1'b0, rs1_i } : 
                                                      (N5)? { 1'b0, 1'b0, 1'b0, rs1_i } : 
                                                      (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N21;
  assign N1 = N24;
  assign N2 = N26;
  assign N3 = N30;
  assign N4 = N33;
  assign N5 = N35;
  assign N6 = N38;
  assign { N67, N66, N65, N64, N63, N62, N61, N60 } = (N0)? data_i : 
                                                      (N1)? data_i : 
                                                      (N2)? { N39, N40, N41, N42, N43, N44, N45, N46 } : 
                                                      (N3)? { 1'b0, 1'b0, 1'b0, rs1_i } : 
                                                      (N4)? { 1'b0, 1'b0, 1'b0, rs1_i } : 
                                                      (N5)? { 1'b0, 1'b0, 1'b0, N47, N48, N49, N50, N51 } : 
                                                      (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign write_data = (N7)? { N67, N66, N65, N64, N63, N62, N61, N60 } : 
                      (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = v_i;
  assign N8 = N85;
  assign write_mask = (N7)? { N59, N58, N57, N56, N55, N54, N53, N52 } : 
                      (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N81, N80, N79 } = (N9)? write_mask[2:0] : 
                             (N10)? write_mask[7:5] : 1'b0;
  assign N9 = N125;
  assign N10 = addr_i[0];
  assign { N84, N83, N82 } = (N9)? write_data[2:0] : 
                             (N10)? write_data[7:5] : 1'b0;
  assign frm_write_mask = (N11)? { N81, N80, N79 } : 
                          (N12)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N78;
  assign N12 = N77;
  assign frm_write_data = (N11)? { N84, N83, N82 } : 
                          (N12)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N93, N92, N91, N90, N89 } = (N13)? write_data[4:0] : 
                                       (N88)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N87;
  assign { N98, N97, N96, N95, N94 } = (N13)? write_mask[4:0] : 
                                       (N88)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign fflags_write_data = (N7)? { N93, N92, N91, N90, N89 } : 
                             (N8)? combined_fflags : 1'b0;
  assign fflags_write_mask = (N7)? { N98, N97, N96, N95, N94 } : 
                             (N8)? combined_fflags : 1'b0;
  assign { N134, N133, N132, N131, N130, N129, N128, N127 } = (N14)? { 1'b0, 1'b0, 1'b0, fflags_r } : 
                                                              (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, frm_o } : 
                                                              (N16)? { frm_o, fflags_r } : 
                                                              (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = N120;
  assign N15 = N122;
  assign N16 = N123;
  assign N17 = N126;
  assign N135 = (N14)? 1'b1 : 
                (N15)? 1'b1 : 
                (N16)? 1'b1 : 
                (N17)? 1'b0 : 1'b0;
  assign data_o = (N18)? { N134, N133, N132, N131, N130, N129, N128, N127 } : 
                  (N118)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = N117;
  assign data_v_o = (N18)? N135 : 
                    (N118)? 1'b0 : 1'b0;
  assign N21 = ~N20;
  assign N24 = ~N23;
  assign N26 = ~N25;
  assign N27 = ~funct3_i[2];
  assign N30 = ~N29;
  assign N33 = ~N32;
  assign N36 = ~funct3_i[1];
  assign N37 = ~funct3_i[0];
  assign N39 = ~data_i[7];
  assign N40 = ~data_i[6];
  assign N41 = ~data_i[5];
  assign N42 = ~data_i[4];
  assign N43 = ~data_i[3];
  assign N44 = ~data_i[2];
  assign N45 = ~data_i[1];
  assign N46 = ~data_i[0];
  assign N47 = ~rs1_i[4];
  assign N48 = ~rs1_i[3];
  assign N49 = ~rs1_i[2];
  assign N50 = ~rs1_i[1];
  assign N51 = ~rs1_i[0];
  assign N78 = ~N77;
  assign filtered_fflags[4] = fflags_v_i[0] & fflags_i[4];
  assign filtered_fflags[3] = fflags_v_i[0] & fflags_i[3];
  assign filtered_fflags[2] = fflags_v_i[0] & fflags_i[2];
  assign filtered_fflags[1] = fflags_v_i[0] & fflags_i[1];
  assign filtered_fflags[0] = fflags_v_i[0] & fflags_i[0];
  assign filtered_fflags[9] = fflags_v_i[1] & fflags_i[9];
  assign filtered_fflags[8] = fflags_v_i[1] & fflags_i[8];
  assign filtered_fflags[7] = fflags_v_i[1] & fflags_i[7];
  assign filtered_fflags[6] = fflags_v_i[1] & fflags_i[6];
  assign filtered_fflags[5] = fflags_v_i[1] & fflags_i[5];
  assign combined_fflags[4] = filtered_fflags[4] | filtered_fflags[9];
  assign combined_fflags[3] = filtered_fflags[3] | filtered_fflags[8];
  assign combined_fflags[2] = filtered_fflags[2] | filtered_fflags[7];
  assign combined_fflags[1] = filtered_fflags[1] | filtered_fflags[6];
  assign combined_fflags[0] = filtered_fflags[0] | filtered_fflags[5];
  assign N85 = ~v_i;
  assign N88 = ~N87;
  assign N99 = ~addr_i[11];
  assign N100 = ~addr_i[10];
  assign N101 = ~addr_i[9];
  assign N102 = ~addr_i[8];
  assign N103 = ~addr_i[7];
  assign N104 = ~addr_i[6];
  assign N105 = ~addr_i[5];
  assign N106 = ~addr_i[4];
  assign N107 = ~addr_i[3];
  assign N108 = ~addr_i[2];
  assign N118 = ~N117;
  assign N120 = ~N119;
  assign N122 = ~N121;
  assign N124 = ~addr_i[1];
  assign N125 = ~addr_i[0];

  always @(posedge clk_i) begin
    if(reset_i) begin
      fflags_r_4_sv2v_reg <= 1'b0;
    end else if(fflags_write_mask[4]) begin
      fflags_r_4_sv2v_reg <= fflags_write_data[4];
    end 
    if(reset_i) begin
      fflags_r_3_sv2v_reg <= 1'b0;
    end else if(fflags_write_mask[3]) begin
      fflags_r_3_sv2v_reg <= fflags_write_data[3];
    end 
    if(reset_i) begin
      fflags_r_2_sv2v_reg <= 1'b0;
    end else if(fflags_write_mask[2]) begin
      fflags_r_2_sv2v_reg <= fflags_write_data[2];
    end 
    if(reset_i) begin
      fflags_r_1_sv2v_reg <= 1'b0;
    end else if(fflags_write_mask[1]) begin
      fflags_r_1_sv2v_reg <= fflags_write_data[1];
    end 
    if(reset_i) begin
      fflags_r_0_sv2v_reg <= 1'b0;
    end else if(fflags_write_mask[0]) begin
      fflags_r_0_sv2v_reg <= fflags_write_data[0];
    end 
    if(reset_i) begin
      frm_o_2_sv2v_reg <= 1'b0;
    end else if(frm_write_mask[2]) begin
      frm_o_2_sv2v_reg <= frm_write_data[2];
    end 
    if(reset_i) begin
      frm_o_1_sv2v_reg <= 1'b0;
    end else if(frm_write_mask[1]) begin
      frm_o_1_sv2v_reg <= frm_write_data[1];
    end 
    if(reset_i) begin
      frm_o_0_sv2v_reg <= 1'b0;
    end else if(frm_write_mask[0]) begin
      frm_o_0_sv2v_reg <= frm_write_data[0];
    end 
  end


endmodule



module mcsr_pc_width_p22_credit_counter_width_p6_cfg_pod_width_p7
(
  clk_i,
  reset_i,
  remote_interrupt_set_i,
  remote_interrupt_clear_i,
  we_i,
  addr_i,
  funct3_i,
  data_i,
  rs1_i,
  data_o,
  cfg_pod_reset_val_i,
  cfg_pod_r_o,
  instr_executed_i,
  interrupt_entered_i,
  mret_called_i,
  npc_r_i,
  mepc_r_o,
  credit_limit_o,
  mstatus_r_o_mpie_,
  mstatus_r_o_mie_,
  mip_r_o_trace_,
  mip_r_o_remote_,
  mie_r_o_trace_,
  mie_r_o_remote_
);

  input [11:0] addr_i;
  input [2:0] funct3_i;
  input [31:0] data_i;
  input [4:0] rs1_i;
  output [31:0] data_o;
  input [6:0] cfg_pod_reset_val_i;
  output [6:0] cfg_pod_r_o;
  input [21:0] npc_r_i;
  output [21:0] mepc_r_o;
  output [5:0] credit_limit_o;
  input clk_i;
  input reset_i;
  input remote_interrupt_set_i;
  input remote_interrupt_clear_i;
  input we_i;
  input instr_executed_i;
  input interrupt_entered_i;
  input mret_called_i;
  output mstatus_r_o_mpie_;
  output mstatus_r_o_mie_;
  output mip_r_o_trace_;
  output mip_r_o_remote_;
  output mie_r_o_trace_;
  output mie_r_o_remote_;
  wire [31:0] data_o;
  wire [6:0] cfg_pod_r_o;
  wire [21:0] mepc_r_o,mepc_n;
  wire [5:0] credit_limit_o;
  wire mstatus_r_o_mpie_,mstatus_r_o_mie_,mip_r_o_trace_,mip_r_o_remote_,
  mie_r_o_trace_,mie_r_o_remote_,N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,mstatus_n_mpie_,mstatus_n_mie_,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,mip_n_remote_,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,
  N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,
  N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,
  N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,
  N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
  N219,N2,N3,N7,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,
  N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,
  N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,
  N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,
  N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,
  N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,
  N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,
  N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,
  N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,
  N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
  N489;
  reg cfg_pod_r_o_6_sv2v_reg,cfg_pod_r_o_5_sv2v_reg,cfg_pod_r_o_4_sv2v_reg,
  cfg_pod_r_o_3_sv2v_reg,cfg_pod_r_o_2_sv2v_reg,cfg_pod_r_o_1_sv2v_reg,
  cfg_pod_r_o_0_sv2v_reg,credit_limit_o_5_sv2v_reg,credit_limit_o_4_sv2v_reg,credit_limit_o_3_sv2v_reg,
  credit_limit_o_2_sv2v_reg,credit_limit_o_1_sv2v_reg,credit_limit_o_0_sv2v_reg,
  mstatus_r_o_mpie__sv2v_reg,mstatus_r_o_mie__sv2v_reg,mie_r_o_trace__sv2v_reg,
  mie_r_o_remote__sv2v_reg,mip_r_o_trace__sv2v_reg,mip_r_o_remote__sv2v_reg,
  mepc_r_o_21_sv2v_reg,mepc_r_o_20_sv2v_reg,mepc_r_o_19_sv2v_reg,mepc_r_o_18_sv2v_reg,
  mepc_r_o_17_sv2v_reg,mepc_r_o_16_sv2v_reg,mepc_r_o_15_sv2v_reg,mepc_r_o_14_sv2v_reg,
  mepc_r_o_13_sv2v_reg,mepc_r_o_12_sv2v_reg,mepc_r_o_11_sv2v_reg,mepc_r_o_10_sv2v_reg,
  mepc_r_o_9_sv2v_reg,mepc_r_o_8_sv2v_reg,mepc_r_o_7_sv2v_reg,mepc_r_o_6_sv2v_reg,
  mepc_r_o_5_sv2v_reg,mepc_r_o_4_sv2v_reg,mepc_r_o_3_sv2v_reg,mepc_r_o_2_sv2v_reg,
  mepc_r_o_1_sv2v_reg,mepc_r_o_0_sv2v_reg;
  assign cfg_pod_r_o[6] = cfg_pod_r_o_6_sv2v_reg;
  assign cfg_pod_r_o[5] = cfg_pod_r_o_5_sv2v_reg;
  assign cfg_pod_r_o[4] = cfg_pod_r_o_4_sv2v_reg;
  assign cfg_pod_r_o[3] = cfg_pod_r_o_3_sv2v_reg;
  assign cfg_pod_r_o[2] = cfg_pod_r_o_2_sv2v_reg;
  assign cfg_pod_r_o[1] = cfg_pod_r_o_1_sv2v_reg;
  assign cfg_pod_r_o[0] = cfg_pod_r_o_0_sv2v_reg;
  assign credit_limit_o[5] = credit_limit_o_5_sv2v_reg;
  assign credit_limit_o[4] = credit_limit_o_4_sv2v_reg;
  assign credit_limit_o[3] = credit_limit_o_3_sv2v_reg;
  assign credit_limit_o[2] = credit_limit_o_2_sv2v_reg;
  assign credit_limit_o[1] = credit_limit_o_1_sv2v_reg;
  assign credit_limit_o[0] = credit_limit_o_0_sv2v_reg;
  assign mstatus_r_o_mpie_ = mstatus_r_o_mpie__sv2v_reg;
  assign mstatus_r_o_mie_ = mstatus_r_o_mie__sv2v_reg;
  assign mie_r_o_trace_ = mie_r_o_trace__sv2v_reg;
  assign mie_r_o_remote_ = mie_r_o_remote__sv2v_reg;
  assign mip_r_o_trace_ = mip_r_o_trace__sv2v_reg;
  assign mip_r_o_remote_ = mip_r_o_remote__sv2v_reg;
  assign mepc_r_o[21] = mepc_r_o_21_sv2v_reg;
  assign mepc_r_o[20] = mepc_r_o_20_sv2v_reg;
  assign mepc_r_o[19] = mepc_r_o_19_sv2v_reg;
  assign mepc_r_o[18] = mepc_r_o_18_sv2v_reg;
  assign mepc_r_o[17] = mepc_r_o_17_sv2v_reg;
  assign mepc_r_o[16] = mepc_r_o_16_sv2v_reg;
  assign mepc_r_o[15] = mepc_r_o_15_sv2v_reg;
  assign mepc_r_o[14] = mepc_r_o_14_sv2v_reg;
  assign mepc_r_o[13] = mepc_r_o_13_sv2v_reg;
  assign mepc_r_o[12] = mepc_r_o_12_sv2v_reg;
  assign mepc_r_o[11] = mepc_r_o_11_sv2v_reg;
  assign mepc_r_o[10] = mepc_r_o_10_sv2v_reg;
  assign mepc_r_o[9] = mepc_r_o_9_sv2v_reg;
  assign mepc_r_o[8] = mepc_r_o_8_sv2v_reg;
  assign mepc_r_o[7] = mepc_r_o_7_sv2v_reg;
  assign mepc_r_o[6] = mepc_r_o_6_sv2v_reg;
  assign mepc_r_o[5] = mepc_r_o_5_sv2v_reg;
  assign mepc_r_o[4] = mepc_r_o_4_sv2v_reg;
  assign mepc_r_o[3] = mepc_r_o_3_sv2v_reg;
  assign mepc_r_o[2] = mepc_r_o_2_sv2v_reg;
  assign mepc_r_o[1] = mepc_r_o_1_sv2v_reg;
  assign mepc_r_o[0] = mepc_r_o_0_sv2v_reg;
  assign data_o[24] = 1'b0;
  assign data_o[25] = 1'b0;
  assign data_o[26] = 1'b0;
  assign data_o[27] = 1'b0;
  assign data_o[28] = 1'b0;
  assign data_o[29] = 1'b0;
  assign data_o[30] = 1'b0;
  assign data_o[31] = 1'b0;
  assign N46 = funct3_i[2] | funct3_i[1];
  assign N47 = N46 | N446;
  assign N49 = funct3_i[2] | N87;
  assign N50 = N49 | funct3_i[0];
  assign N52 = N49 | N446;
  assign N54 = N83 | funct3_i[1];
  assign N55 = N54 | N446;
  assign N57 = N83 | N87;
  assign N58 = N57 | funct3_i[0];
  assign N60 = funct3_i[2] & funct3_i[1];
  assign N61 = N60 & funct3_i[0];
  assign N74 = funct3_i[1] | N446;
  assign N84 = N87 | funct3_i[0];
  assign N86 = funct3_i[1] & funct3_i[0];
  assign N88 = N87 & N446;
  assign N153 = addr_i[9] & addr_i[8];
  assign N154 = N150 & N151;
  assign N155 = N153 & N154;
  assign N156 = N155 & N152;
  assign N158 = N428 & N429;
  assign N159 = N432 & N433;
  assign N160 = N450 & N463;
  assign N161 = N158 & N159;
  assign N162 = N160 & N483;
  assign N163 = N161 & N162;
  assign N164 = addr_i[7] | addr_i[6];
  assign N165 = N182 | N164;
  assign N166 = N165 | N169;
  assign N168 = addr_i[5] | N463;
  assign N169 = N168 | addr_i[0];
  assign N170 = N185 | N169;
  assign N172 = N177 | N483;
  assign N173 = N185 | N172;
  assign N175 = N428 | N429;
  assign N176 = N432 | N433;
  assign N177 = addr_i[5] | addr_i[2];
  assign N178 = N175 | N176;
  assign N179 = N177 | addr_i[0];
  assign N180 = N178 | N179;
  assign N182 = addr_i[11] | addr_i[10];
  assign N183 = addr_i[7] | N433;
  assign N184 = N450 | addr_i[2];
  assign N185 = N182 | N183;
  assign N186 = N184 | addr_i[0];
  assign N187 = N185 | N186;
  assign N220 = reset_i | mret_called_i;
  assign N428 = ~addr_i[11];
  assign N429 = ~addr_i[10];
  assign N430 = ~addr_i[9];
  assign N431 = ~addr_i[8];
  assign N432 = ~addr_i[7];
  assign N433 = ~addr_i[6];
  assign N434 = N429 | N428;
  assign N435 = N430 | N434;
  assign N436 = N431 | N435;
  assign N437 = N432 | N436;
  assign N438 = N433 | N437;
  assign N439 = addr_i[5] | N438;
  assign N440 = addr_i[4] | N439;
  assign N441 = addr_i[3] | N440;
  assign N442 = addr_i[2] | N441;
  assign N443 = addr_i[1] | N442;
  assign N444 = addr_i[0] | N443;
  assign N445 = ~N444;
  assign N446 = ~funct3_i[0];
  assign N447 = funct3_i[1] | funct3_i[2];
  assign N448 = N446 | N447;
  assign N449 = ~N448;
  assign N450 = ~addr_i[5];
  assign N451 = addr_i[10] | addr_i[11];
  assign N452 = N430 | N451;
  assign N453 = N431 | N452;
  assign N454 = addr_i[7] | N453;
  assign N455 = N433 | N454;
  assign N456 = N450 | N455;
  assign N457 = addr_i[4] | N456;
  assign N458 = addr_i[3] | N457;
  assign N459 = addr_i[2] | N458;
  assign N460 = addr_i[1] | N459;
  assign N461 = addr_i[0] | N460;
  assign N462 = ~N461;
  assign N463 = ~addr_i[2];
  assign N464 = addr_i[5] | N455;
  assign N465 = addr_i[4] | N464;
  assign N466 = addr_i[3] | N465;
  assign N467 = N463 | N466;
  assign N468 = addr_i[1] | N467;
  assign N469 = addr_i[0] | N468;
  assign N470 = ~N469;
  assign N471 = addr_i[6] | N454;
  assign N472 = addr_i[5] | N471;
  assign N473 = addr_i[4] | N472;
  assign N474 = addr_i[3] | N473;
  assign N475 = N463 | N474;
  assign N476 = addr_i[1] | N475;
  assign N477 = addr_i[0] | N476;
  assign N478 = ~N477;
  assign N479 = addr_i[2] | N474;
  assign N480 = addr_i[1] | N479;
  assign N481 = addr_i[0] | N480;
  assign N482 = ~N481;
  assign N483 = ~addr_i[0];
  assign N484 = addr_i[2] | N466;
  assign N485 = addr_i[1] | N484;
  assign N486 = N483 | N485;
  assign N487 = ~N486;
  assign N32 = (N0)? 1'b1 : 
               (N41)? 1'b1 : 
               (N31)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign { N39, N38, N37, N36, N35, N34, N33 } = (N0)? cfg_pod_reset_val_i : 
                                                 (N41)? data_i[6:0] : 1'b0;
  assign N63 = (N1)? 1'b1 : 
               (N62)? mstatus_r_o_mpie_ : 1'b0;
  assign N1 = data_i[7];
  assign N64 = (N1)? 1'b0 : 
               (N62)? mstatus_r_o_mpie_ : 1'b0;
  assign N66 = (N4)? data_i[3] : 
               (N5)? 1'b1 : 
               (N6)? 1'b0 : 
               (N8)? rs1_i[3] : 
               (N9)? 1'b1 : 
               (N10)? 1'b0 : 1'b0;
  assign N4 = N48;
  assign N5 = N51;
  assign N6 = N53;
  assign N8 = N56;
  assign N9 = N59;
  assign N10 = N61;
  assign N67 = (N4)? data_i[7] : 
               (N5)? N63 : 
               (N6)? N64 : 
               (N8)? mstatus_r_o_mpie_ : 
               (N9)? mstatus_r_o_mpie_ : 
               (N10)? mstatus_r_o_mpie_ : 
               (N11)? mstatus_r_o_mpie_ : 1'b0;
  assign N11 = N88;
  assign mstatus_n_mie_ = (N12)? mstatus_r_o_mpie_ : 
                          (N69)? 1'b0 : 
                          (N71)? N66 : 1'b0;
  assign N12 = mret_called_i;
  assign mstatus_n_mpie_ = (N13)? mstatus_r_o_mie_ : 
                           (N7)? N67 : 
                           (N3)? mstatus_r_o_mpie_ : 1'b0;
  assign N13 = interrupt_entered_i;
  assign { N78, N77 } = (N14)? data_i[17:16] : 
                        (N15)? { 1'b1, 1'b1 } : 
                        (N16)? { 1'b0, 1'b0 } : 1'b0;
  assign N14 = N75;
  assign N15 = N85;
  assign N16 = N86;
  assign N90 = (N17)? 1'b1 : 
               (N89)? mip_r_o_trace_ : 1'b0;
  assign N17 = data_i[17];
  assign N91 = (N17)? 1'b0 : 
               (N89)? mip_r_o_trace_ : 1'b0;
  assign N92 = (N14)? data_i[17] : 
               (N15)? N90 : 
               (N16)? N91 : 
               (N11)? mip_r_o_trace_ : 1'b0;
  assign N93 = (N18)? N92 : 
               (N19)? mip_r_o_trace_ : 1'b0;
  assign N18 = N83;
  assign N19 = funct3_i[2];
  assign N94 = (N20)? 1'b1 : 
               (N99)? N93 : 
               (N82)? mip_r_o_trace_ : 1'b0;
  assign N20 = N79;
  assign mip_n_remote_ = (N21)? 1'b1 : 
                         (N101)? 1'b0 : 
                         (N104)? N77 : 1'b0;
  assign N21 = remote_interrupt_set_i;
  assign { N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127 } = (N14)? { data_i[23:18], data_i[15:2] } : 
                                                                                                                                      (N15)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                      (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign mepc_n = (N13)? npc_r_i : 
                  (N148)? { N146, N145, N144, N143, N142, N141, N78, N77, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127 } : 1'b0;
  assign { N213, N212, N202, N201, N200, N199, N198, N197, N196, N195 } = (N22)? { 1'b0, 1'b0, mstatus_r_o_mpie_, 1'b0, 1'b0, 1'b0, mstatus_r_o_mie_, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N23)? { mie_r_o_trace_, mie_r_o_remote_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N24)? { mip_r_o_trace_, mip_r_o_remote_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N25)? { mepc_r_o[15:14], mepc_r_o[5:0], 1'b0, 1'b0 } : 
                                                                          (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, credit_limit_o } : 
                                                                          (N27)? { 1'b0, 1'b0, 1'b0, cfg_pod_r_o } : 
                                                                          (N194)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = N163;
  assign N23 = N167;
  assign N24 = N171;
  assign N25 = N174;
  assign N26 = N181;
  assign N27 = N188;
  assign { N219, N218, N217, N216, N215, N214, N211, N210, N209, N208, N207, N206, N205, N204 } = (N25)? { mepc_r_o[21:16], mepc_r_o[13:6] } : 
                                                                                                  (N203)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_o[23:0] = (N28)? { N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N202, N201, N200, N199, N198, N197, N196, N195 } : 
                        (N157)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N28 = N156;
  assign N29 = N488 & N449;
  assign N488 = we_i & N462;
  assign N30 = N29 | reset_i;
  assign N31 = ~N30;
  assign N40 = ~reset_i;
  assign N41 = N29 & N40;
  assign N42 = we_i & N482;
  assign N43 = interrupt_entered_i | mret_called_i;
  assign N44 = N42 | N43;
  assign N45 = ~N44;
  assign N48 = ~N47;
  assign N51 = ~N50;
  assign N53 = ~N52;
  assign N56 = ~N55;
  assign N59 = ~N58;
  assign N62 = ~data_i[7];
  assign N65 = ~rs1_i[3];
  assign N68 = ~mret_called_i;
  assign N69 = interrupt_entered_i & N68;
  assign N70 = N68 & N147;
  assign N71 = N42 & N70;
  assign N72 = we_i & N478;
  assign N73 = ~N72;
  assign N75 = ~N74;
  assign N76 = ~data_i[16];
  assign N79 = instr_executed_i & mie_r_o_trace_;
  assign N80 = we_i & N470;
  assign N81 = N80 | N79;
  assign N82 = ~N81;
  assign N83 = ~funct3_i[2];
  assign N85 = ~N84;
  assign N87 = ~funct3_i[1];
  assign N89 = ~data_i[17];
  assign N95 = remote_interrupt_clear_i | remote_interrupt_set_i;
  assign N96 = N80 | N95;
  assign N97 = ~N96;
  assign N98 = ~N79;
  assign N99 = N80 & N98;
  assign N100 = ~remote_interrupt_set_i;
  assign N101 = remote_interrupt_clear_i & N100;
  assign N102 = ~remote_interrupt_clear_i;
  assign N103 = N100 & N102;
  assign N104 = N80 & N103;
  assign N105 = we_i & N487;
  assign N106 = N105 | interrupt_entered_i;
  assign N107 = ~N106;
  assign N108 = ~data_i[2];
  assign N109 = ~data_i[3];
  assign N110 = ~data_i[4];
  assign N111 = ~data_i[5];
  assign N112 = ~data_i[6];
  assign N113 = ~data_i[8];
  assign N114 = ~data_i[9];
  assign N115 = ~data_i[10];
  assign N116 = ~data_i[11];
  assign N117 = ~data_i[12];
  assign N118 = ~data_i[13];
  assign N119 = ~data_i[14];
  assign N120 = ~data_i[15];
  assign N121 = ~data_i[18];
  assign N122 = ~data_i[19];
  assign N123 = ~data_i[20];
  assign N124 = ~data_i[21];
  assign N125 = ~data_i[22];
  assign N126 = ~data_i[23];
  assign N147 = ~interrupt_entered_i;
  assign N148 = N105 & N147;
  assign N149 = N489 & N449;
  assign N489 = we_i & N445;
  assign N150 = ~addr_i[4];
  assign N151 = ~addr_i[3];
  assign N152 = ~addr_i[1];
  assign N157 = ~N156;
  assign N167 = ~N166;
  assign N171 = ~N170;
  assign N174 = ~N173;
  assign N181 = ~N180;
  assign N188 = ~N187;
  assign N189 = N167 | N163;
  assign N190 = N171 | N189;
  assign N191 = N174 | N190;
  assign N192 = N181 | N191;
  assign N193 = N188 | N192;
  assign N194 = ~N193;
  assign N203 = N173;
  assign N2 = N42 | interrupt_entered_i;
  assign N3 = ~N2;
  assign N7 = N42 & N147;
  assign N221 = N51 & N71;
  assign N222 = N109 & N221;
  assign N223 = N53 & N71;
  assign N224 = N109 & N223;
  assign N225 = N222 | N224;
  assign N226 = N59 & N71;
  assign N227 = N65 & N226;
  assign N228 = N225 | N227;
  assign N229 = N61 & N71;
  assign N230 = N65 & N229;
  assign N231 = N228 | N230;
  assign N232 = N88 & N71;
  assign N233 = N231 | N232;
  assign N234 = N233 | N45;
  assign N235 = ~N234;
  assign N236 = N83 & N72;
  assign N237 = N85 & N236;
  assign N238 = N89 & N237;
  assign N239 = N86 & N236;
  assign N240 = N89 & N239;
  assign N241 = N238 | N240;
  assign N242 = N88 & N236;
  assign N243 = N241 | N242;
  assign N244 = funct3_i[2] & N72;
  assign N245 = N243 | N244;
  assign N246 = N245 | N73;
  assign N247 = ~N246;
  assign N248 = N76 & N237;
  assign N249 = N76 & N239;
  assign N250 = N248 | N249;
  assign N251 = N250 | N242;
  assign N252 = N251 | N244;
  assign N253 = N252 | N73;
  assign N254 = ~N253;
  assign N255 = N83 & N104;
  assign N256 = N88 & N255;
  assign N257 = funct3_i[2] & N104;
  assign N258 = N256 | N257;
  assign N259 = ~N258;
  assign N260 = N85 & N255;
  assign N261 = N76 & N260;
  assign N262 = N86 & N255;
  assign N263 = N76 & N262;
  assign N264 = N261 | N263;
  assign N265 = N264 | N256;
  assign N266 = N265 | N257;
  assign N267 = N266 | N97;
  assign N268 = ~N267;
  assign N269 = N83 & N148;
  assign N270 = N85 & N269;
  assign N271 = N126 & N270;
  assign N272 = N86 & N269;
  assign N273 = N126 & N272;
  assign N274 = N271 | N273;
  assign N275 = N88 & N269;
  assign N276 = N274 | N275;
  assign N277 = funct3_i[2] & N148;
  assign N278 = N276 | N277;
  assign N279 = N278 | N107;
  assign N280 = ~N279;
  assign N281 = N125 & N270;
  assign N282 = N125 & N272;
  assign N283 = N281 | N282;
  assign N284 = N283 | N275;
  assign N285 = N284 | N277;
  assign N286 = N285 | N107;
  assign N287 = ~N286;
  assign N288 = N124 & N270;
  assign N289 = N124 & N272;
  assign N290 = N288 | N289;
  assign N291 = N290 | N275;
  assign N292 = N291 | N277;
  assign N293 = N292 | N107;
  assign N294 = ~N293;
  assign N295 = N123 & N270;
  assign N296 = N123 & N272;
  assign N297 = N295 | N296;
  assign N298 = N297 | N275;
  assign N299 = N298 | N277;
  assign N300 = N299 | N107;
  assign N301 = ~N300;
  assign N302 = N122 & N270;
  assign N303 = N122 & N272;
  assign N304 = N302 | N303;
  assign N305 = N304 | N275;
  assign N306 = N305 | N277;
  assign N307 = N306 | N107;
  assign N308 = ~N307;
  assign N309 = N121 & N270;
  assign N310 = N121 & N272;
  assign N311 = N309 | N310;
  assign N312 = N311 | N275;
  assign N313 = N312 | N277;
  assign N314 = N313 | N107;
  assign N315 = ~N314;
  assign N316 = N89 & N270;
  assign N317 = N89 & N272;
  assign N318 = N316 | N317;
  assign N319 = N318 | N275;
  assign N320 = N319 | N277;
  assign N321 = N320 | N107;
  assign N322 = ~N321;
  assign N323 = N76 & N270;
  assign N324 = N76 & N272;
  assign N325 = N323 | N324;
  assign N326 = N325 | N275;
  assign N327 = N326 | N277;
  assign N328 = N327 | N107;
  assign N329 = ~N328;
  assign N330 = N120 & N270;
  assign N331 = N120 & N272;
  assign N332 = N330 | N331;
  assign N333 = N332 | N275;
  assign N334 = N333 | N277;
  assign N335 = N334 | N107;
  assign N336 = ~N335;
  assign N337 = N119 & N270;
  assign N338 = N119 & N272;
  assign N339 = N337 | N338;
  assign N340 = N339 | N275;
  assign N341 = N340 | N277;
  assign N342 = N341 | N107;
  assign N343 = ~N342;
  assign N344 = N118 & N270;
  assign N345 = N118 & N272;
  assign N346 = N344 | N345;
  assign N347 = N346 | N275;
  assign N348 = N347 | N277;
  assign N349 = N348 | N107;
  assign N350 = ~N349;
  assign N351 = N117 & N270;
  assign N352 = N117 & N272;
  assign N353 = N351 | N352;
  assign N354 = N353 | N275;
  assign N355 = N354 | N277;
  assign N356 = N355 | N107;
  assign N357 = ~N356;
  assign N358 = N116 & N270;
  assign N359 = N116 & N272;
  assign N360 = N358 | N359;
  assign N361 = N360 | N275;
  assign N362 = N361 | N277;
  assign N363 = N362 | N107;
  assign N364 = ~N363;
  assign N365 = N115 & N270;
  assign N366 = N115 & N272;
  assign N367 = N365 | N366;
  assign N368 = N367 | N275;
  assign N369 = N368 | N277;
  assign N370 = N369 | N107;
  assign N371 = ~N370;
  assign N372 = N114 & N270;
  assign N373 = N114 & N272;
  assign N374 = N372 | N373;
  assign N375 = N374 | N275;
  assign N376 = N375 | N277;
  assign N377 = N376 | N107;
  assign N378 = ~N377;
  assign N379 = N113 & N270;
  assign N380 = N113 & N272;
  assign N381 = N379 | N380;
  assign N382 = N381 | N275;
  assign N383 = N382 | N277;
  assign N384 = N383 | N107;
  assign N385 = ~N384;
  assign N386 = N62 & N270;
  assign N387 = N62 & N272;
  assign N388 = N386 | N387;
  assign N389 = N388 | N275;
  assign N390 = N389 | N277;
  assign N391 = N390 | N107;
  assign N392 = ~N391;
  assign N393 = N112 & N270;
  assign N394 = N112 & N272;
  assign N395 = N393 | N394;
  assign N396 = N395 | N275;
  assign N397 = N396 | N277;
  assign N398 = N397 | N107;
  assign N399 = ~N398;
  assign N400 = N111 & N270;
  assign N401 = N111 & N272;
  assign N402 = N400 | N401;
  assign N403 = N402 | N275;
  assign N404 = N403 | N277;
  assign N405 = N404 | N107;
  assign N406 = ~N405;
  assign N407 = N110 & N270;
  assign N408 = N110 & N272;
  assign N409 = N407 | N408;
  assign N410 = N409 | N275;
  assign N411 = N410 | N277;
  assign N412 = N411 | N107;
  assign N413 = ~N412;
  assign N414 = N109 & N270;
  assign N415 = N109 & N272;
  assign N416 = N414 | N415;
  assign N417 = N416 | N275;
  assign N418 = N417 | N277;
  assign N419 = N418 | N107;
  assign N420 = ~N419;
  assign N421 = N108 & N270;
  assign N422 = N108 & N272;
  assign N423 = N421 | N422;
  assign N424 = N423 | N275;
  assign N425 = N424 | N277;
  assign N426 = N425 | N107;
  assign N427 = ~N426;

  always @(posedge clk_i) begin
    if(N32) begin
      cfg_pod_r_o_6_sv2v_reg <= N39;
      cfg_pod_r_o_5_sv2v_reg <= N38;
      cfg_pod_r_o_4_sv2v_reg <= N37;
      cfg_pod_r_o_3_sv2v_reg <= N36;
      cfg_pod_r_o_2_sv2v_reg <= N35;
      cfg_pod_r_o_1_sv2v_reg <= N34;
      cfg_pod_r_o_0_sv2v_reg <= N33;
    end 
    if(reset_i) begin
      credit_limit_o_5_sv2v_reg <= 1'b1;
      credit_limit_o_4_sv2v_reg <= 1'b0;
      credit_limit_o_3_sv2v_reg <= 1'b0;
      credit_limit_o_2_sv2v_reg <= 1'b0;
      credit_limit_o_1_sv2v_reg <= 1'b0;
      credit_limit_o_0_sv2v_reg <= 1'b0;
    end else if(N149) begin
      credit_limit_o_5_sv2v_reg <= data_i[5];
      credit_limit_o_4_sv2v_reg <= data_i[4];
      credit_limit_o_3_sv2v_reg <= data_i[3];
      credit_limit_o_2_sv2v_reg <= data_i[2];
      credit_limit_o_1_sv2v_reg <= data_i[1];
      credit_limit_o_0_sv2v_reg <= data_i[0];
    end 
    if(N220) begin
      mstatus_r_o_mpie__sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      mstatus_r_o_mpie__sv2v_reg <= mstatus_n_mpie_;
    end 
    if(reset_i) begin
      mstatus_r_o_mie__sv2v_reg <= 1'b0;
    end else if(N235) begin
      mstatus_r_o_mie__sv2v_reg <= mstatus_n_mie_;
    end 
    if(reset_i) begin
      mie_r_o_trace__sv2v_reg <= 1'b0;
    end else if(N247) begin
      mie_r_o_trace__sv2v_reg <= N78;
    end 
    if(reset_i) begin
      mie_r_o_remote__sv2v_reg <= 1'b0;
    end else if(N254) begin
      mie_r_o_remote__sv2v_reg <= N77;
    end 
    if(reset_i) begin
      mip_r_o_trace__sv2v_reg <= 1'b0;
    end else if(N259) begin
      mip_r_o_trace__sv2v_reg <= N94;
    end 
    if(reset_i) begin
      mip_r_o_remote__sv2v_reg <= 1'b0;
    end else if(N268) begin
      mip_r_o_remote__sv2v_reg <= mip_n_remote_;
    end 
    if(reset_i) begin
      mepc_r_o_21_sv2v_reg <= 1'b0;
    end else if(N280) begin
      mepc_r_o_21_sv2v_reg <= mepc_n[21];
    end 
    if(reset_i) begin
      mepc_r_o_20_sv2v_reg <= 1'b0;
    end else if(N287) begin
      mepc_r_o_20_sv2v_reg <= mepc_n[20];
    end 
    if(reset_i) begin
      mepc_r_o_19_sv2v_reg <= 1'b0;
    end else if(N294) begin
      mepc_r_o_19_sv2v_reg <= mepc_n[19];
    end 
    if(reset_i) begin
      mepc_r_o_18_sv2v_reg <= 1'b0;
    end else if(N301) begin
      mepc_r_o_18_sv2v_reg <= mepc_n[18];
    end 
    if(reset_i) begin
      mepc_r_o_17_sv2v_reg <= 1'b0;
    end else if(N308) begin
      mepc_r_o_17_sv2v_reg <= mepc_n[17];
    end 
    if(reset_i) begin
      mepc_r_o_16_sv2v_reg <= 1'b0;
    end else if(N315) begin
      mepc_r_o_16_sv2v_reg <= mepc_n[16];
    end 
    if(reset_i) begin
      mepc_r_o_15_sv2v_reg <= 1'b0;
    end else if(N322) begin
      mepc_r_o_15_sv2v_reg <= mepc_n[15];
    end 
    if(reset_i) begin
      mepc_r_o_14_sv2v_reg <= 1'b0;
    end else if(N329) begin
      mepc_r_o_14_sv2v_reg <= mepc_n[14];
    end 
    if(reset_i) begin
      mepc_r_o_13_sv2v_reg <= 1'b0;
    end else if(N336) begin
      mepc_r_o_13_sv2v_reg <= mepc_n[13];
    end 
    if(reset_i) begin
      mepc_r_o_12_sv2v_reg <= 1'b0;
    end else if(N343) begin
      mepc_r_o_12_sv2v_reg <= mepc_n[12];
    end 
    if(reset_i) begin
      mepc_r_o_11_sv2v_reg <= 1'b0;
    end else if(N350) begin
      mepc_r_o_11_sv2v_reg <= mepc_n[11];
    end 
    if(reset_i) begin
      mepc_r_o_10_sv2v_reg <= 1'b0;
    end else if(N357) begin
      mepc_r_o_10_sv2v_reg <= mepc_n[10];
    end 
    if(reset_i) begin
      mepc_r_o_9_sv2v_reg <= 1'b0;
    end else if(N364) begin
      mepc_r_o_9_sv2v_reg <= mepc_n[9];
    end 
    if(reset_i) begin
      mepc_r_o_8_sv2v_reg <= 1'b0;
    end else if(N371) begin
      mepc_r_o_8_sv2v_reg <= mepc_n[8];
    end 
    if(reset_i) begin
      mepc_r_o_7_sv2v_reg <= 1'b0;
    end else if(N378) begin
      mepc_r_o_7_sv2v_reg <= mepc_n[7];
    end 
    if(reset_i) begin
      mepc_r_o_6_sv2v_reg <= 1'b0;
    end else if(N385) begin
      mepc_r_o_6_sv2v_reg <= mepc_n[6];
    end 
    if(reset_i) begin
      mepc_r_o_5_sv2v_reg <= 1'b0;
    end else if(N392) begin
      mepc_r_o_5_sv2v_reg <= mepc_n[5];
    end 
    if(reset_i) begin
      mepc_r_o_4_sv2v_reg <= 1'b0;
    end else if(N399) begin
      mepc_r_o_4_sv2v_reg <= mepc_n[4];
    end 
    if(reset_i) begin
      mepc_r_o_3_sv2v_reg <= 1'b0;
    end else if(N406) begin
      mepc_r_o_3_sv2v_reg <= mepc_n[3];
    end 
    if(reset_i) begin
      mepc_r_o_2_sv2v_reg <= 1'b0;
    end else if(N413) begin
      mepc_r_o_2_sv2v_reg <= mepc_n[2];
    end 
    if(reset_i) begin
      mepc_r_o_1_sv2v_reg <= 1'b0;
    end else if(N420) begin
      mepc_r_o_1_sv2v_reg <= mepc_n[1];
    end 
    if(reset_i) begin
      mepc_r_o_0_sv2v_reg <= 1'b0;
    end else if(N427) begin
      mepc_r_o_0_sv2v_reg <= mepc_n[0];
    end 
  end


endmodule



module bsg_mux_width_p33_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [65:0] data_i;
  input [0:0] sel_i;
  output [32:0] data_o;
  wire [32:0] data_o;
  wire N0,N1;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[65] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[64] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[63] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[62] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[61] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[60] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[59] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[58] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[57] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[56] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[55] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[54] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[53] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[52] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[51] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[50] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[49] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[48] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[47] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[46] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[45] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[44] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[43] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[42] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[41] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[40] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[39] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[38] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[37] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[36] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[35] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[34] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[33] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module recFNToRawFN_expWidth8_sigWidth24
(
  in,
  isNaN,
  isInf,
  isZero,
  sign,
  sExp,
  sig
);

  input [32:0] in;
  output [9:0] sExp;
  output [24:0] sig;
  output isNaN;
  output isInf;
  output isZero;
  output sign;
  wire [9:0] sExp;
  wire [24:0] sig;
  wire isNaN,isInf,isZero,sign,in_32_,sExp_8_,sExp_7_,sExp_6_,sExp_5_,sExp_4_,sExp_3_,
  sExp_2_,sExp_1_,sExp_0_,sig_22_,sig_21_,sig_20_,sig_19_,sig_18_,sig_17_,sig_16_,
  sig_15_,sig_14_,sig_13_,sig_12_,sig_11_,sig_10_,sig_9_,sig_8_,sig_7_,sig_6_,
  sig_5_,sig_4_,sig_3_,sig_2_,sig_1_,sig_0_,N0,N1,N2,N4;
  assign sig[24] = 1'b0;
  assign sExp[9] = 1'b0;
  assign in_32_ = in[32];
  assign sign = in_32_;
  assign sExp_8_ = in[31];
  assign sExp[8] = sExp_8_;
  assign sExp_7_ = in[30];
  assign sExp[7] = sExp_7_;
  assign sExp_6_ = in[29];
  assign sExp[6] = sExp_6_;
  assign sExp_5_ = in[28];
  assign sExp[5] = sExp_5_;
  assign sExp_4_ = in[27];
  assign sExp[4] = sExp_4_;
  assign sExp_3_ = in[26];
  assign sExp[3] = sExp_3_;
  assign sExp_2_ = in[25];
  assign sExp[2] = sExp_2_;
  assign sExp_1_ = in[24];
  assign sExp[1] = sExp_1_;
  assign sExp_0_ = in[23];
  assign sExp[0] = sExp_0_;
  assign sig_22_ = in[22];
  assign sig[22] = sig_22_;
  assign sig_21_ = in[21];
  assign sig[21] = sig_21_;
  assign sig_20_ = in[20];
  assign sig[20] = sig_20_;
  assign sig_19_ = in[19];
  assign sig[19] = sig_19_;
  assign sig_18_ = in[18];
  assign sig[18] = sig_18_;
  assign sig_17_ = in[17];
  assign sig[17] = sig_17_;
  assign sig_16_ = in[16];
  assign sig[16] = sig_16_;
  assign sig_15_ = in[15];
  assign sig[15] = sig_15_;
  assign sig_14_ = in[14];
  assign sig[14] = sig_14_;
  assign sig_13_ = in[13];
  assign sig[13] = sig_13_;
  assign sig_12_ = in[12];
  assign sig[12] = sig_12_;
  assign sig_11_ = in[11];
  assign sig[11] = sig_11_;
  assign sig_10_ = in[10];
  assign sig[10] = sig_10_;
  assign sig_9_ = in[9];
  assign sig[9] = sig_9_;
  assign sig_8_ = in[8];
  assign sig[8] = sig_8_;
  assign sig_7_ = in[7];
  assign sig[7] = sig_7_;
  assign sig_6_ = in[6];
  assign sig[6] = sig_6_;
  assign sig_5_ = in[5];
  assign sig[5] = sig_5_;
  assign sig_4_ = in[4];
  assign sig[4] = sig_4_;
  assign sig_3_ = in[3];
  assign sig[3] = sig_3_;
  assign sig_2_ = in[2];
  assign sig[2] = sig_2_;
  assign sig_1_ = in[1];
  assign sig[1] = sig_1_;
  assign sig_0_ = in[0];
  assign sig[0] = sig_0_;
  assign N0 = sExp_7_ & sExp_8_;
  assign N1 = sExp_7_ | sExp_8_;
  assign N2 = sExp_6_ | N1;
  assign isZero = ~N2;
  assign isNaN = N0 & sExp_6_;
  assign isInf = N0 & N4;
  assign N4 = ~sExp_6_;
  assign sig[23] = ~isZero;

endmodule



module recFNToFN_expWidth8_sigWidth24
(
  in,
  out
);

  input [32:0] in;
  output [31:0] out;
  wire [31:0] out;
  wire N0,N1,isNaN,isInf,isZero,N2,isSubnormal,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,sv2v_dc_1;
  wire [9:0] sExp;
  wire [24:0] sig;
  wire [4:0] denormShiftDist;

  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN
  (
    .in(in),
    .isNaN(isNaN),
    .isInf(isInf),
    .isZero(isZero),
    .sign(out[31]),
    .sExp(sExp),
    .sig(sig)
  );

  assign N2 = sExp[5:0] <= 1'b1;
  assign N56 = ~sExp[7];
  assign N57 = sExp[8] | sExp[9];
  assign N58 = N56 | N57;
  assign N59 = sExp[6] | N58;
  assign N60 = ~N59;
  assign N61 = sExp[8] | sExp[9];
  assign N62 = sExp[7] | N61;
  assign N63 = ~N62;
  assign denormShiftDist = 1'b1 - sExp[4:0];
  assign { sv2v_dc_1, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31 } = sig[24:1] >> denormShiftDist;
  assign { N11, N10, N9, N8, N7, N6, N5, N4 } = sExp[7:0] - { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign { N19, N18, N17, N16, N15, N14, N13, N12 } = { N11, N10, N9, N8, N7, N6, N5, N4 } + 1'b1;
  assign { N27, N26, N25, N24, N23, N22, N21, N20 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N1)? { N19, N18, N17, N16, N15, N14, N13, N12 } : 1'b0;
  assign N0 = isSubnormal;
  assign N1 = N3;
  assign out[22:0] = (N0)? { N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31 } : 
                     (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N30)? sig[22:0] : 1'b0;
  assign isSubnormal = N64 | N63;
  assign N64 = N60 & N2;
  assign N3 = ~isSubnormal;
  assign N28 = isNaN | isInf;
  assign out[30] = N27 | N28;
  assign out[29] = N26 | N28;
  assign out[28] = N25 | N28;
  assign out[27] = N24 | N28;
  assign out[26] = N23 | N28;
  assign out[25] = N22 | N28;
  assign out[24] = N21 | N28;
  assign out[23] = N20 | N28;
  assign N29 = isInf | isSubnormal;
  assign N30 = ~N29;
  assign N54 = ~isSubnormal;
  assign N55 = isInf & N54;

endmodule



module bsg_mux_width_p32_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [95:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[31] = (N2)? data_i[31] : 
                      (N3)? data_i[63] : 
                      (N4)? data_i[95] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[30] = (N2)? data_i[30] : 
                      (N3)? data_i[62] : 
                      (N4)? data_i[94] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N3)? data_i[61] : 
                      (N4)? data_i[93] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N3)? data_i[60] : 
                      (N4)? data_i[92] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N3)? data_i[59] : 
                      (N4)? data_i[91] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N3)? data_i[58] : 
                      (N4)? data_i[90] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N3)? data_i[57] : 
                      (N4)? data_i[89] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N3)? data_i[56] : 
                      (N4)? data_i[88] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N3)? data_i[55] : 
                      (N4)? data_i[87] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N3)? data_i[54] : 
                      (N4)? data_i[86] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N3)? data_i[53] : 
                      (N4)? data_i[85] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N3)? data_i[52] : 
                      (N4)? data_i[84] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N3)? data_i[51] : 
                      (N4)? data_i[83] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N3)? data_i[50] : 
                      (N4)? data_i[82] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N3)? data_i[49] : 
                      (N4)? data_i[81] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N3)? data_i[48] : 
                      (N4)? data_i[80] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N3)? data_i[47] : 
                      (N4)? data_i[79] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N3)? data_i[46] : 
                      (N4)? data_i[78] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N3)? data_i[45] : 
                      (N4)? data_i[77] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N3)? data_i[44] : 
                      (N4)? data_i[76] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N3)? data_i[43] : 
                      (N4)? data_i[75] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N3)? data_i[42] : 
                      (N4)? data_i[74] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N3)? data_i[41] : 
                     (N4)? data_i[73] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N3)? data_i[40] : 
                     (N4)? data_i[72] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N3)? data_i[39] : 
                     (N4)? data_i[71] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N3)? data_i[38] : 
                     (N4)? data_i[70] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N3)? data_i[37] : 
                     (N4)? data_i[69] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N3)? data_i[36] : 
                     (N4)? data_i[68] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[35] : 
                     (N4)? data_i[67] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[34] : 
                     (N4)? data_i[66] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[33] : 
                     (N4)? data_i[65] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[32] : 
                     (N4)? data_i[64] : 1'b0;

endmodule



module bsg_dff_reset_width_p225
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [224:0] data_i;
  output [224:0] data_o;
  input clk_i;
  input reset_i;
  wire [224:0] data_o;
  reg data_o_224_sv2v_reg,data_o_223_sv2v_reg,data_o_222_sv2v_reg,data_o_221_sv2v_reg,
  data_o_220_sv2v_reg,data_o_219_sv2v_reg,data_o_218_sv2v_reg,data_o_217_sv2v_reg,
  data_o_216_sv2v_reg,data_o_215_sv2v_reg,data_o_214_sv2v_reg,data_o_213_sv2v_reg,
  data_o_212_sv2v_reg,data_o_211_sv2v_reg,data_o_210_sv2v_reg,data_o_209_sv2v_reg,
  data_o_208_sv2v_reg,data_o_207_sv2v_reg,data_o_206_sv2v_reg,data_o_205_sv2v_reg,
  data_o_204_sv2v_reg,data_o_203_sv2v_reg,data_o_202_sv2v_reg,data_o_201_sv2v_reg,
  data_o_200_sv2v_reg,data_o_199_sv2v_reg,data_o_198_sv2v_reg,data_o_197_sv2v_reg,
  data_o_196_sv2v_reg,data_o_195_sv2v_reg,data_o_194_sv2v_reg,data_o_193_sv2v_reg,
  data_o_192_sv2v_reg,data_o_191_sv2v_reg,data_o_190_sv2v_reg,data_o_189_sv2v_reg,
  data_o_188_sv2v_reg,data_o_187_sv2v_reg,data_o_186_sv2v_reg,data_o_185_sv2v_reg,
  data_o_184_sv2v_reg,data_o_183_sv2v_reg,data_o_182_sv2v_reg,data_o_181_sv2v_reg,
  data_o_180_sv2v_reg,data_o_179_sv2v_reg,data_o_178_sv2v_reg,data_o_177_sv2v_reg,
  data_o_176_sv2v_reg,data_o_175_sv2v_reg,data_o_174_sv2v_reg,data_o_173_sv2v_reg,
  data_o_172_sv2v_reg,data_o_171_sv2v_reg,data_o_170_sv2v_reg,data_o_169_sv2v_reg,
  data_o_168_sv2v_reg,data_o_167_sv2v_reg,data_o_166_sv2v_reg,data_o_165_sv2v_reg,
  data_o_164_sv2v_reg,data_o_163_sv2v_reg,data_o_162_sv2v_reg,data_o_161_sv2v_reg,
  data_o_160_sv2v_reg,data_o_159_sv2v_reg,data_o_158_sv2v_reg,data_o_157_sv2v_reg,
  data_o_156_sv2v_reg,data_o_155_sv2v_reg,data_o_154_sv2v_reg,data_o_153_sv2v_reg,
  data_o_152_sv2v_reg,data_o_151_sv2v_reg,data_o_150_sv2v_reg,data_o_149_sv2v_reg,
  data_o_148_sv2v_reg,data_o_147_sv2v_reg,data_o_146_sv2v_reg,data_o_145_sv2v_reg,
  data_o_144_sv2v_reg,data_o_143_sv2v_reg,data_o_142_sv2v_reg,data_o_141_sv2v_reg,
  data_o_140_sv2v_reg,data_o_139_sv2v_reg,data_o_138_sv2v_reg,data_o_137_sv2v_reg,
  data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,data_o_133_sv2v_reg,
  data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,data_o_129_sv2v_reg,
  data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,data_o_125_sv2v_reg,
  data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,data_o_121_sv2v_reg,
  data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,data_o_117_sv2v_reg,
  data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,data_o_113_sv2v_reg,
  data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,data_o_109_sv2v_reg,
  data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,data_o_105_sv2v_reg,
  data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,data_o_101_sv2v_reg,
  data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,data_o_97_sv2v_reg,
  data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,data_o_93_sv2v_reg,
  data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,data_o_89_sv2v_reg,
  data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,data_o_85_sv2v_reg,
  data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,
  data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,
  data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,
  data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_224_sv2v_reg <= 1'b0;
      data_o_223_sv2v_reg <= 1'b0;
      data_o_222_sv2v_reg <= 1'b0;
      data_o_221_sv2v_reg <= 1'b0;
      data_o_220_sv2v_reg <= 1'b0;
      data_o_219_sv2v_reg <= 1'b0;
      data_o_218_sv2v_reg <= 1'b0;
      data_o_217_sv2v_reg <= 1'b0;
      data_o_216_sv2v_reg <= 1'b0;
      data_o_215_sv2v_reg <= 1'b0;
      data_o_214_sv2v_reg <= 1'b0;
      data_o_213_sv2v_reg <= 1'b0;
      data_o_212_sv2v_reg <= 1'b0;
      data_o_211_sv2v_reg <= 1'b0;
      data_o_210_sv2v_reg <= 1'b0;
      data_o_209_sv2v_reg <= 1'b0;
      data_o_208_sv2v_reg <= 1'b0;
      data_o_207_sv2v_reg <= 1'b0;
      data_o_206_sv2v_reg <= 1'b0;
      data_o_205_sv2v_reg <= 1'b0;
      data_o_204_sv2v_reg <= 1'b0;
      data_o_203_sv2v_reg <= 1'b0;
      data_o_202_sv2v_reg <= 1'b0;
      data_o_201_sv2v_reg <= 1'b0;
      data_o_200_sv2v_reg <= 1'b0;
      data_o_199_sv2v_reg <= 1'b0;
      data_o_198_sv2v_reg <= 1'b0;
      data_o_197_sv2v_reg <= 1'b0;
      data_o_196_sv2v_reg <= 1'b0;
      data_o_195_sv2v_reg <= 1'b0;
      data_o_194_sv2v_reg <= 1'b0;
      data_o_193_sv2v_reg <= 1'b0;
      data_o_192_sv2v_reg <= 1'b0;
      data_o_191_sv2v_reg <= 1'b0;
      data_o_190_sv2v_reg <= 1'b0;
      data_o_189_sv2v_reg <= 1'b0;
      data_o_188_sv2v_reg <= 1'b0;
      data_o_187_sv2v_reg <= 1'b0;
      data_o_186_sv2v_reg <= 1'b0;
      data_o_185_sv2v_reg <= 1'b0;
      data_o_184_sv2v_reg <= 1'b0;
      data_o_183_sv2v_reg <= 1'b0;
      data_o_182_sv2v_reg <= 1'b0;
      data_o_181_sv2v_reg <= 1'b0;
      data_o_180_sv2v_reg <= 1'b0;
      data_o_179_sv2v_reg <= 1'b0;
      data_o_178_sv2v_reg <= 1'b0;
      data_o_177_sv2v_reg <= 1'b0;
      data_o_176_sv2v_reg <= 1'b0;
      data_o_175_sv2v_reg <= 1'b0;
      data_o_174_sv2v_reg <= 1'b0;
      data_o_173_sv2v_reg <= 1'b0;
      data_o_172_sv2v_reg <= 1'b0;
      data_o_171_sv2v_reg <= 1'b0;
      data_o_170_sv2v_reg <= 1'b0;
      data_o_169_sv2v_reg <= 1'b0;
      data_o_168_sv2v_reg <= 1'b0;
      data_o_167_sv2v_reg <= 1'b0;
      data_o_166_sv2v_reg <= 1'b0;
      data_o_165_sv2v_reg <= 1'b0;
      data_o_164_sv2v_reg <= 1'b0;
      data_o_163_sv2v_reg <= 1'b0;
      data_o_162_sv2v_reg <= 1'b0;
      data_o_161_sv2v_reg <= 1'b0;
      data_o_160_sv2v_reg <= 1'b0;
      data_o_159_sv2v_reg <= 1'b0;
      data_o_158_sv2v_reg <= 1'b0;
      data_o_157_sv2v_reg <= 1'b0;
      data_o_156_sv2v_reg <= 1'b0;
      data_o_155_sv2v_reg <= 1'b0;
      data_o_154_sv2v_reg <= 1'b0;
      data_o_153_sv2v_reg <= 1'b0;
      data_o_152_sv2v_reg <= 1'b0;
      data_o_151_sv2v_reg <= 1'b0;
      data_o_150_sv2v_reg <= 1'b0;
      data_o_149_sv2v_reg <= 1'b0;
      data_o_148_sv2v_reg <= 1'b0;
      data_o_147_sv2v_reg <= 1'b0;
      data_o_146_sv2v_reg <= 1'b0;
      data_o_145_sv2v_reg <= 1'b0;
      data_o_144_sv2v_reg <= 1'b0;
      data_o_143_sv2v_reg <= 1'b0;
      data_o_142_sv2v_reg <= 1'b0;
      data_o_141_sv2v_reg <= 1'b0;
      data_o_140_sv2v_reg <= 1'b0;
      data_o_139_sv2v_reg <= 1'b0;
      data_o_138_sv2v_reg <= 1'b0;
      data_o_137_sv2v_reg <= 1'b0;
      data_o_136_sv2v_reg <= 1'b0;
      data_o_135_sv2v_reg <= 1'b0;
      data_o_134_sv2v_reg <= 1'b0;
      data_o_133_sv2v_reg <= 1'b0;
      data_o_132_sv2v_reg <= 1'b0;
      data_o_131_sv2v_reg <= 1'b0;
      data_o_130_sv2v_reg <= 1'b0;
      data_o_129_sv2v_reg <= 1'b0;
      data_o_128_sv2v_reg <= 1'b0;
      data_o_127_sv2v_reg <= 1'b0;
      data_o_126_sv2v_reg <= 1'b0;
      data_o_125_sv2v_reg <= 1'b0;
      data_o_124_sv2v_reg <= 1'b0;
      data_o_123_sv2v_reg <= 1'b0;
      data_o_122_sv2v_reg <= 1'b0;
      data_o_121_sv2v_reg <= 1'b0;
      data_o_120_sv2v_reg <= 1'b0;
      data_o_119_sv2v_reg <= 1'b0;
      data_o_118_sv2v_reg <= 1'b0;
      data_o_117_sv2v_reg <= 1'b0;
      data_o_116_sv2v_reg <= 1'b0;
      data_o_115_sv2v_reg <= 1'b0;
      data_o_114_sv2v_reg <= 1'b0;
      data_o_113_sv2v_reg <= 1'b0;
      data_o_112_sv2v_reg <= 1'b0;
      data_o_111_sv2v_reg <= 1'b0;
      data_o_110_sv2v_reg <= 1'b0;
      data_o_109_sv2v_reg <= 1'b0;
      data_o_108_sv2v_reg <= 1'b0;
      data_o_107_sv2v_reg <= 1'b0;
      data_o_106_sv2v_reg <= 1'b0;
      data_o_105_sv2v_reg <= 1'b0;
      data_o_104_sv2v_reg <= 1'b0;
      data_o_103_sv2v_reg <= 1'b0;
      data_o_102_sv2v_reg <= 1'b0;
      data_o_101_sv2v_reg <= 1'b0;
      data_o_100_sv2v_reg <= 1'b0;
      data_o_99_sv2v_reg <= 1'b0;
      data_o_98_sv2v_reg <= 1'b0;
      data_o_97_sv2v_reg <= 1'b0;
      data_o_96_sv2v_reg <= 1'b0;
      data_o_95_sv2v_reg <= 1'b0;
      data_o_94_sv2v_reg <= 1'b0;
      data_o_93_sv2v_reg <= 1'b0;
      data_o_92_sv2v_reg <= 1'b0;
      data_o_91_sv2v_reg <= 1'b0;
      data_o_90_sv2v_reg <= 1'b0;
      data_o_89_sv2v_reg <= 1'b0;
      data_o_88_sv2v_reg <= 1'b0;
      data_o_87_sv2v_reg <= 1'b0;
      data_o_86_sv2v_reg <= 1'b0;
      data_o_85_sv2v_reg <= 1'b0;
      data_o_84_sv2v_reg <= 1'b0;
      data_o_83_sv2v_reg <= 1'b0;
      data_o_82_sv2v_reg <= 1'b0;
      data_o_81_sv2v_reg <= 1'b0;
      data_o_80_sv2v_reg <= 1'b0;
      data_o_79_sv2v_reg <= 1'b0;
      data_o_78_sv2v_reg <= 1'b0;
      data_o_77_sv2v_reg <= 1'b0;
      data_o_76_sv2v_reg <= 1'b0;
      data_o_75_sv2v_reg <= 1'b0;
      data_o_74_sv2v_reg <= 1'b0;
      data_o_73_sv2v_reg <= 1'b0;
      data_o_72_sv2v_reg <= 1'b0;
      data_o_71_sv2v_reg <= 1'b0;
      data_o_70_sv2v_reg <= 1'b0;
      data_o_69_sv2v_reg <= 1'b0;
      data_o_68_sv2v_reg <= 1'b0;
      data_o_67_sv2v_reg <= 1'b0;
      data_o_66_sv2v_reg <= 1'b0;
      data_o_65_sv2v_reg <= 1'b0;
      data_o_64_sv2v_reg <= 1'b0;
      data_o_63_sv2v_reg <= 1'b0;
      data_o_62_sv2v_reg <= 1'b0;
      data_o_61_sv2v_reg <= 1'b0;
      data_o_60_sv2v_reg <= 1'b0;
      data_o_59_sv2v_reg <= 1'b0;
      data_o_58_sv2v_reg <= 1'b0;
      data_o_57_sv2v_reg <= 1'b0;
      data_o_56_sv2v_reg <= 1'b0;
      data_o_55_sv2v_reg <= 1'b0;
      data_o_54_sv2v_reg <= 1'b0;
      data_o_53_sv2v_reg <= 1'b0;
      data_o_52_sv2v_reg <= 1'b0;
      data_o_51_sv2v_reg <= 1'b0;
      data_o_50_sv2v_reg <= 1'b0;
      data_o_49_sv2v_reg <= 1'b0;
      data_o_48_sv2v_reg <= 1'b0;
      data_o_47_sv2v_reg <= 1'b0;
      data_o_46_sv2v_reg <= 1'b0;
      data_o_45_sv2v_reg <= 1'b0;
      data_o_44_sv2v_reg <= 1'b0;
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_224_sv2v_reg <= data_i[224];
      data_o_223_sv2v_reg <= data_i[223];
      data_o_222_sv2v_reg <= data_i[222];
      data_o_221_sv2v_reg <= data_i[221];
      data_o_220_sv2v_reg <= data_i[220];
      data_o_219_sv2v_reg <= data_i[219];
      data_o_218_sv2v_reg <= data_i[218];
      data_o_217_sv2v_reg <= data_i[217];
      data_o_216_sv2v_reg <= data_i[216];
      data_o_215_sv2v_reg <= data_i[215];
      data_o_214_sv2v_reg <= data_i[214];
      data_o_213_sv2v_reg <= data_i[213];
      data_o_212_sv2v_reg <= data_i[212];
      data_o_211_sv2v_reg <= data_i[211];
      data_o_210_sv2v_reg <= data_i[210];
      data_o_209_sv2v_reg <= data_i[209];
      data_o_208_sv2v_reg <= data_i[208];
      data_o_207_sv2v_reg <= data_i[207];
      data_o_206_sv2v_reg <= data_i[206];
      data_o_205_sv2v_reg <= data_i[205];
      data_o_204_sv2v_reg <= data_i[204];
      data_o_203_sv2v_reg <= data_i[203];
      data_o_202_sv2v_reg <= data_i[202];
      data_o_201_sv2v_reg <= data_i[201];
      data_o_200_sv2v_reg <= data_i[200];
      data_o_199_sv2v_reg <= data_i[199];
      data_o_198_sv2v_reg <= data_i[198];
      data_o_197_sv2v_reg <= data_i[197];
      data_o_196_sv2v_reg <= data_i[196];
      data_o_195_sv2v_reg <= data_i[195];
      data_o_194_sv2v_reg <= data_i[194];
      data_o_193_sv2v_reg <= data_i[193];
      data_o_192_sv2v_reg <= data_i[192];
      data_o_191_sv2v_reg <= data_i[191];
      data_o_190_sv2v_reg <= data_i[190];
      data_o_189_sv2v_reg <= data_i[189];
      data_o_188_sv2v_reg <= data_i[188];
      data_o_187_sv2v_reg <= data_i[187];
      data_o_186_sv2v_reg <= data_i[186];
      data_o_185_sv2v_reg <= data_i[185];
      data_o_184_sv2v_reg <= data_i[184];
      data_o_183_sv2v_reg <= data_i[183];
      data_o_182_sv2v_reg <= data_i[182];
      data_o_181_sv2v_reg <= data_i[181];
      data_o_180_sv2v_reg <= data_i[180];
      data_o_179_sv2v_reg <= data_i[179];
      data_o_178_sv2v_reg <= data_i[178];
      data_o_177_sv2v_reg <= data_i[177];
      data_o_176_sv2v_reg <= data_i[176];
      data_o_175_sv2v_reg <= data_i[175];
      data_o_174_sv2v_reg <= data_i[174];
      data_o_173_sv2v_reg <= data_i[173];
      data_o_172_sv2v_reg <= data_i[172];
      data_o_171_sv2v_reg <= data_i[171];
      data_o_170_sv2v_reg <= data_i[170];
      data_o_169_sv2v_reg <= data_i[169];
      data_o_168_sv2v_reg <= data_i[168];
      data_o_167_sv2v_reg <= data_i[167];
      data_o_166_sv2v_reg <= data_i[166];
      data_o_165_sv2v_reg <= data_i[165];
      data_o_164_sv2v_reg <= data_i[164];
      data_o_163_sv2v_reg <= data_i[163];
      data_o_162_sv2v_reg <= data_i[162];
      data_o_161_sv2v_reg <= data_i[161];
      data_o_160_sv2v_reg <= data_i[160];
      data_o_159_sv2v_reg <= data_i[159];
      data_o_158_sv2v_reg <= data_i[158];
      data_o_157_sv2v_reg <= data_i[157];
      data_o_156_sv2v_reg <= data_i[156];
      data_o_155_sv2v_reg <= data_i[155];
      data_o_154_sv2v_reg <= data_i[154];
      data_o_153_sv2v_reg <= data_i[153];
      data_o_152_sv2v_reg <= data_i[152];
      data_o_151_sv2v_reg <= data_i[151];
      data_o_150_sv2v_reg <= data_i[150];
      data_o_149_sv2v_reg <= data_i[149];
      data_o_148_sv2v_reg <= data_i[148];
      data_o_147_sv2v_reg <= data_i[147];
      data_o_146_sv2v_reg <= data_i[146];
      data_o_145_sv2v_reg <= data_i[145];
      data_o_144_sv2v_reg <= data_i[144];
      data_o_143_sv2v_reg <= data_i[143];
      data_o_142_sv2v_reg <= data_i[142];
      data_o_141_sv2v_reg <= data_i[141];
      data_o_140_sv2v_reg <= data_i[140];
      data_o_139_sv2v_reg <= data_i[139];
      data_o_138_sv2v_reg <= data_i[138];
      data_o_137_sv2v_reg <= data_i[137];
      data_o_136_sv2v_reg <= data_i[136];
      data_o_135_sv2v_reg <= data_i[135];
      data_o_134_sv2v_reg <= data_i[134];
      data_o_133_sv2v_reg <= data_i[133];
      data_o_132_sv2v_reg <= data_i[132];
      data_o_131_sv2v_reg <= data_i[131];
      data_o_130_sv2v_reg <= data_i[130];
      data_o_129_sv2v_reg <= data_i[129];
      data_o_128_sv2v_reg <= data_i[128];
      data_o_127_sv2v_reg <= data_i[127];
      data_o_126_sv2v_reg <= data_i[126];
      data_o_125_sv2v_reg <= data_i[125];
      data_o_124_sv2v_reg <= data_i[124];
      data_o_123_sv2v_reg <= data_i[123];
      data_o_122_sv2v_reg <= data_i[122];
      data_o_121_sv2v_reg <= data_i[121];
      data_o_120_sv2v_reg <= data_i[120];
      data_o_119_sv2v_reg <= data_i[119];
      data_o_118_sv2v_reg <= data_i[118];
      data_o_117_sv2v_reg <= data_i[117];
      data_o_116_sv2v_reg <= data_i[116];
      data_o_115_sv2v_reg <= data_i[115];
      data_o_114_sv2v_reg <= data_i[114];
      data_o_113_sv2v_reg <= data_i[113];
      data_o_112_sv2v_reg <= data_i[112];
      data_o_111_sv2v_reg <= data_i[111];
      data_o_110_sv2v_reg <= data_i[110];
      data_o_109_sv2v_reg <= data_i[109];
      data_o_108_sv2v_reg <= data_i[108];
      data_o_107_sv2v_reg <= data_i[107];
      data_o_106_sv2v_reg <= data_i[106];
      data_o_105_sv2v_reg <= data_i[105];
      data_o_104_sv2v_reg <= data_i[104];
      data_o_103_sv2v_reg <= data_i[103];
      data_o_102_sv2v_reg <= data_i[102];
      data_o_101_sv2v_reg <= data_i[101];
      data_o_100_sv2v_reg <= data_i[100];
      data_o_99_sv2v_reg <= data_i[99];
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module alu_pc_width_p22
(
  rs1_i,
  rs2_i,
  pc_plus4_i,
  op_i,
  result_o,
  jalr_addr_o,
  jump_now_o
);

  input [31:0] rs1_i;
  input [31:0] rs2_i;
  input [31:0] pc_plus4_i;
  input [31:0] op_i;
  output [31:0] result_o;
  output [21:0] jalr_addr_o;
  output jump_now_o;
  wire [31:0] result_o,op2,adder_input,shr_out,shl_out,xor_out,and_out,or_out;
  wire [21:0] jalr_addr_o;
  wire jump_now_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,is_imm_op,N26,sub_not_add,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  carry,sign_ex_or_zero,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,
  N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,
  N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,
  N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
  N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,
  N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,
  N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,
  N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,
  N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,rs1_eq_rs2,
  rs1_lt_rs2_unsigned,rs1_lt_rs2_signed,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,sv2v_dc_1;
  wire [4:0] sh_amount;
  wire [32:0] sum;
  assign { sv2v_dc_1, shr_out } = $signed({ sign_ex_or_zero, rs1_i }) >>> sh_amount;
  assign shl_out = rs1_i << sh_amount;
  assign N94 = op_i[6] | N329;
  assign N95 = N94 | N99;
  assign N96 = N95 | N212;
  assign N98 = op_i[6] | op_i[5];
  assign N99 = N319 | op_i[3];
  assign N100 = N98 | N99;
  assign N101 = N100 | N212;
  assign N103 = N303 & N127;
  assign N104 = N103 & N141;
  assign N105 = N104 & N203;
  assign N106 = N150 & N197;
  assign N107 = N106 & op_i[0];
  assign N109 = N313 & N127;
  assign N110 = N109 & N141;
  assign N111 = N110 & N203;
  assign N112 = N150 & N133;
  assign N113 = N112 & op_i[0];
  assign N115 = N313 & N137;
  assign N116 = N115 & N141;
  assign N117 = N116 & N203;
  assign N118 = N150 & N146;
  assign N119 = N118 & op_i[0];
  assign N121 = N306 & N127;
  assign N122 = N121 & N141;
  assign N123 = N122 & N203;
  assign N124 = N159 & N197;
  assign N125 = N124 & op_i[0];
  assign N127 = N302 & N328;
  assign N128 = N309 & N127;
  assign N129 = N128 & N141;
  assign N130 = N129 & N203;
  assign N131 = op_i[13] & N302;
  assign N132 = N131 & N190;
  assign N133 = N132 & N195;
  assign N134 = N159 & N133;
  assign N135 = N134 & op_i[0];
  assign N137 = op_i[12] & N328;
  assign N138 = N329 & op_i[4];
  assign N139 = N294 & N333;
  assign N140 = N309 & N137;
  assign N141 = N138 & N139;
  assign N142 = N140 & N141;
  assign N143 = N142 & N203;
  assign N144 = op_i[13] & op_i[12];
  assign N145 = N144 & N190;
  assign N146 = N145 & N195;
  assign N147 = N159 & N146;
  assign N148 = N147 & op_i[0];
  assign N150 = N158 & N193;
  assign N151 = N150 & N171;
  assign N152 = N151 & op_i[0];
  assign N153 = N150 & N175;
  assign N154 = N153 & op_i[0];
  assign N157 = N179 & N156;
  assign N158 = N157 & N186;
  assign N159 = N158 & N168;
  assign N160 = N159 & N171;
  assign N161 = N160 & op_i[0];
  assign N162 = N159 & N175;
  assign N163 = N162 & op_i[0];
  assign N165 = N184 & op_i[14];
  assign N166 = N301 & op_i[12];
  assign N167 = N328 & N329;
  assign N168 = N187 & N165;
  assign N169 = N166 & N167;
  assign N170 = N192 & N168;
  assign N171 = N169 & N195;
  assign N172 = N170 & N171;
  assign N173 = N172 & op_i[0];
  assign N174 = N166 & N190;
  assign N175 = N174 & N195;
  assign N176 = N170 & N175;
  assign N177 = N176 & op_i[0];
  assign N185 = N179 & op_i[30];
  assign N186 = N180 & N181;
  assign N187 = N182 & N183;
  assign N188 = N184 & N312;
  assign N189 = N301 & N302;
  assign N190 = N328 & op_i[5];
  assign N191 = op_i[4] & N294;
  assign N192 = N185 & N186;
  assign N193 = N187 & N188;
  assign N194 = N189 & N190;
  assign N195 = N191 & N297;
  assign N196 = N192 & N193;
  assign N197 = N194 & N195;
  assign N198 = N196 & N197;
  assign N199 = N198 & op_i[0];
  assign N200 = N302 & op_i[6];
  assign N201 = op_i[5] & N319;
  assign N202 = N294 & op_i[2];
  assign N203 = op_i[1] & op_i[0];
  assign N204 = N303 & N200;
  assign N205 = N201 & N202;
  assign N206 = N204 & N205;
  assign N207 = N206 & N203;
  assign N208 = N328 | N329;
  assign N209 = op_i[4] | N294;
  assign N210 = N333 | N323;
  assign N211 = N208 | N209;
  assign N212 = N210 | N325;
  assign N213 = N211 | N212;
  assign rs1_eq_rs2 = rs1_i == rs2_i;
  assign rs1_lt_rs2_unsigned = rs1_i < rs2_i;
  assign rs1_lt_rs2_signed = $signed(rs1_i) < $signed(rs2_i);
  assign N295 = op_i[6] & op_i[5];
  assign N296 = N319 & N294;
  assign N297 = N333 & op_i[1];
  assign N298 = N295 & N296;
  assign N299 = N298 & N297;
  assign N303 = N312 & N301;
  assign N304 = N303 & N302;
  assign N305 = N303 & op_i[12];
  assign N306 = op_i[14] & N301;
  assign N307 = N306 & N302;
  assign N308 = N306 & op_i[12];
  assign N309 = op_i[14] & op_i[13];
  assign N310 = N309 & N302;
  assign N311 = N309 & op_i[12];
  assign N313 = N312 & op_i[13];
  assign { N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229 } = { op_i[31:12], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } + pc_plus4_i;
  assign { N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261 } = { N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229 } - { 1'b1, 1'b0, 1'b0 };
  assign { N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60 } = { rs1_i[31:31], rs1_i } + { adder_input[31:31], adder_input };
  assign { carry, sum } = { N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60 } + sub_not_add;
  assign op2 = (N0)? { op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:31], op_i[31:20] } : 
               (N1)? rs2_i : 1'b0;
  assign N0 = is_imm_op;
  assign N1 = N26;
  assign adder_input = (N2)? { N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59 } : 
                       (N3)? op2 : 1'b0;
  assign N2 = sub_not_add;
  assign N3 = N27;
  assign sh_amount = (N0)? op_i[24:20] : 
                     (N1)? rs2_i[4:0] : 1'b0;
  assign result_o = (N4)? { op_i[31:12], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                    (N5)? { N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261 } : 
                    (N6)? sum[31:0] : 
                    (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sum[32:32] } : 
                    (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N293 } : 
                    (N9)? xor_out : 
                    (N10)? or_out : 
                    (N11)? and_out : 
                    (N12)? shl_out : 
                    (N13)? shr_out : 
                    (N14)? shr_out : 
                    (N15)? sum[31:0] : 
                    (N16)? pc_plus4_i : 
                    (N17)? pc_plus4_i : 
                    (N228)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = N97;
  assign N5 = N102;
  assign N6 = N108;
  assign N7 = N114;
  assign N8 = N120;
  assign N9 = N126;
  assign N10 = N136;
  assign N11 = N149;
  assign N12 = N155;
  assign N13 = N164;
  assign N14 = N178;
  assign N15 = N199;
  assign N16 = N207;
  assign N17 = N214;
  assign sub_not_add = (N4)? 1'b0 : 
                       (N5)? 1'b0 : 
                       (N6)? 1'b0 : 
                       (N7)? 1'b1 : 
                       (N8)? 1'b1 : 
                       (N9)? 1'b0 : 
                       (N10)? 1'b0 : 
                       (N11)? 1'b0 : 
                       (N12)? 1'b0 : 
                       (N13)? 1'b0 : 
                       (N14)? 1'b0 : 
                       (N15)? 1'b1 : 
                       (N16)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N228)? 1'b0 : 1'b0;
  assign sign_ex_or_zero = (N4)? 1'b0 : 
                           (N5)? 1'b0 : 
                           (N6)? 1'b0 : 
                           (N7)? 1'b0 : 
                           (N8)? 1'b0 : 
                           (N9)? 1'b0 : 
                           (N10)? 1'b0 : 
                           (N11)? 1'b0 : 
                           (N12)? 1'b0 : 
                           (N13)? 1'b0 : 
                           (N14)? rs1_i[31] : 
                           (N15)? 1'b0 : 
                           (N16)? 1'b0 : 
                           (N17)? 1'b0 : 
                           (N228)? 1'b0 : 1'b0;
  assign jalr_addr_o = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N16)? sum[23:2] : 
                       (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N228)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N317 = (N18)? rs1_eq_rs2 : 
                (N19)? N314 : 
                (N20)? rs1_lt_rs2_signed : 
                (N21)? N315 : 
                (N22)? rs1_lt_rs2_unsigned : 
                (N23)? N316 : 
                (N24)? 1'b0 : 1'b0;
  assign N18 = N304;
  assign N19 = N305;
  assign N20 = N307;
  assign N21 = N308;
  assign N22 = N310;
  assign N23 = N311;
  assign N24 = N313;
  assign jump_now_o = (N25)? N317 : 
                      (N300)? 1'b0 : 1'b0;
  assign N25 = N299;
  assign is_imm_op = N327 | N337;
  assign N327 = ~N326;
  assign N326 = N324 | N325;
  assign N324 = N322 | N323;
  assign N322 = N321 | op_i[2];
  assign N321 = N320 | op_i[3];
  assign N320 = N318 | N319;
  assign N318 = op_i[6] | op_i[5];
  assign N319 = ~op_i[4];
  assign N323 = ~op_i[1];
  assign N325 = ~op_i[0];
  assign N337 = ~N336;
  assign N336 = N335 | N325;
  assign N335 = N334 | N323;
  assign N334 = N332 | N333;
  assign N332 = N331 | op_i[3];
  assign N331 = N330 | op_i[4];
  assign N330 = N328 | N329;
  assign N328 = ~op_i[6];
  assign N329 = ~op_i[5];
  assign N333 = ~op_i[2];
  assign N26 = ~is_imm_op;
  assign N27 = ~sub_not_add;
  assign N28 = ~op2[31];
  assign N29 = ~op2[30];
  assign N30 = ~op2[29];
  assign N31 = ~op2[28];
  assign N32 = ~op2[27];
  assign N33 = ~op2[26];
  assign N34 = ~op2[25];
  assign N35 = ~op2[24];
  assign N36 = ~op2[23];
  assign N37 = ~op2[22];
  assign N38 = ~op2[21];
  assign N39 = ~op2[20];
  assign N40 = ~op2[19];
  assign N41 = ~op2[18];
  assign N42 = ~op2[17];
  assign N43 = ~op2[16];
  assign N44 = ~op2[15];
  assign N45 = ~op2[14];
  assign N46 = ~op2[13];
  assign N47 = ~op2[12];
  assign N48 = ~op2[11];
  assign N49 = ~op2[10];
  assign N50 = ~op2[9];
  assign N51 = ~op2[8];
  assign N52 = ~op2[7];
  assign N53 = ~op2[6];
  assign N54 = ~op2[5];
  assign N55 = ~op2[4];
  assign N56 = ~op2[3];
  assign N57 = ~op2[2];
  assign N58 = ~op2[1];
  assign N59 = ~op2[0];
  assign xor_out[31] = rs1_i[31] ^ op2[31];
  assign xor_out[30] = rs1_i[30] ^ op2[30];
  assign xor_out[29] = rs1_i[29] ^ op2[29];
  assign xor_out[28] = rs1_i[28] ^ op2[28];
  assign xor_out[27] = rs1_i[27] ^ op2[27];
  assign xor_out[26] = rs1_i[26] ^ op2[26];
  assign xor_out[25] = rs1_i[25] ^ op2[25];
  assign xor_out[24] = rs1_i[24] ^ op2[24];
  assign xor_out[23] = rs1_i[23] ^ op2[23];
  assign xor_out[22] = rs1_i[22] ^ op2[22];
  assign xor_out[21] = rs1_i[21] ^ op2[21];
  assign xor_out[20] = rs1_i[20] ^ op2[20];
  assign xor_out[19] = rs1_i[19] ^ op2[19];
  assign xor_out[18] = rs1_i[18] ^ op2[18];
  assign xor_out[17] = rs1_i[17] ^ op2[17];
  assign xor_out[16] = rs1_i[16] ^ op2[16];
  assign xor_out[15] = rs1_i[15] ^ op2[15];
  assign xor_out[14] = rs1_i[14] ^ op2[14];
  assign xor_out[13] = rs1_i[13] ^ op2[13];
  assign xor_out[12] = rs1_i[12] ^ op2[12];
  assign xor_out[11] = rs1_i[11] ^ op2[11];
  assign xor_out[10] = rs1_i[10] ^ op2[10];
  assign xor_out[9] = rs1_i[9] ^ op2[9];
  assign xor_out[8] = rs1_i[8] ^ op2[8];
  assign xor_out[7] = rs1_i[7] ^ op2[7];
  assign xor_out[6] = rs1_i[6] ^ op2[6];
  assign xor_out[5] = rs1_i[5] ^ op2[5];
  assign xor_out[4] = rs1_i[4] ^ op2[4];
  assign xor_out[3] = rs1_i[3] ^ op2[3];
  assign xor_out[2] = rs1_i[2] ^ op2[2];
  assign xor_out[1] = rs1_i[1] ^ op2[1];
  assign xor_out[0] = rs1_i[0] ^ op2[0];
  assign and_out[31] = rs1_i[31] & op2[31];
  assign and_out[30] = rs1_i[30] & op2[30];
  assign and_out[29] = rs1_i[29] & op2[29];
  assign and_out[28] = rs1_i[28] & op2[28];
  assign and_out[27] = rs1_i[27] & op2[27];
  assign and_out[26] = rs1_i[26] & op2[26];
  assign and_out[25] = rs1_i[25] & op2[25];
  assign and_out[24] = rs1_i[24] & op2[24];
  assign and_out[23] = rs1_i[23] & op2[23];
  assign and_out[22] = rs1_i[22] & op2[22];
  assign and_out[21] = rs1_i[21] & op2[21];
  assign and_out[20] = rs1_i[20] & op2[20];
  assign and_out[19] = rs1_i[19] & op2[19];
  assign and_out[18] = rs1_i[18] & op2[18];
  assign and_out[17] = rs1_i[17] & op2[17];
  assign and_out[16] = rs1_i[16] & op2[16];
  assign and_out[15] = rs1_i[15] & op2[15];
  assign and_out[14] = rs1_i[14] & op2[14];
  assign and_out[13] = rs1_i[13] & op2[13];
  assign and_out[12] = rs1_i[12] & op2[12];
  assign and_out[11] = rs1_i[11] & op2[11];
  assign and_out[10] = rs1_i[10] & op2[10];
  assign and_out[9] = rs1_i[9] & op2[9];
  assign and_out[8] = rs1_i[8] & op2[8];
  assign and_out[7] = rs1_i[7] & op2[7];
  assign and_out[6] = rs1_i[6] & op2[6];
  assign and_out[5] = rs1_i[5] & op2[5];
  assign and_out[4] = rs1_i[4] & op2[4];
  assign and_out[3] = rs1_i[3] & op2[3];
  assign and_out[2] = rs1_i[2] & op2[2];
  assign and_out[1] = rs1_i[1] & op2[1];
  assign and_out[0] = rs1_i[0] & op2[0];
  assign or_out[31] = rs1_i[31] | op2[31];
  assign or_out[30] = rs1_i[30] | op2[30];
  assign or_out[29] = rs1_i[29] | op2[29];
  assign or_out[28] = rs1_i[28] | op2[28];
  assign or_out[27] = rs1_i[27] | op2[27];
  assign or_out[26] = rs1_i[26] | op2[26];
  assign or_out[25] = rs1_i[25] | op2[25];
  assign or_out[24] = rs1_i[24] | op2[24];
  assign or_out[23] = rs1_i[23] | op2[23];
  assign or_out[22] = rs1_i[22] | op2[22];
  assign or_out[21] = rs1_i[21] | op2[21];
  assign or_out[20] = rs1_i[20] | op2[20];
  assign or_out[19] = rs1_i[19] | op2[19];
  assign or_out[18] = rs1_i[18] | op2[18];
  assign or_out[17] = rs1_i[17] | op2[17];
  assign or_out[16] = rs1_i[16] | op2[16];
  assign or_out[15] = rs1_i[15] | op2[15];
  assign or_out[14] = rs1_i[14] | op2[14];
  assign or_out[13] = rs1_i[13] | op2[13];
  assign or_out[12] = rs1_i[12] | op2[12];
  assign or_out[11] = rs1_i[11] | op2[11];
  assign or_out[10] = rs1_i[10] | op2[10];
  assign or_out[9] = rs1_i[9] | op2[9];
  assign or_out[8] = rs1_i[8] | op2[8];
  assign or_out[7] = rs1_i[7] | op2[7];
  assign or_out[6] = rs1_i[6] | op2[6];
  assign or_out[5] = rs1_i[5] | op2[5];
  assign or_out[4] = rs1_i[4] | op2[4];
  assign or_out[3] = rs1_i[3] | op2[3];
  assign or_out[2] = rs1_i[2] | op2[2];
  assign or_out[1] = rs1_i[1] | op2[1];
  assign or_out[0] = rs1_i[0] | op2[0];
  assign N97 = ~N96;
  assign N102 = ~N101;
  assign N108 = N105 | N107;
  assign N114 = N111 | N113;
  assign N120 = N117 | N119;
  assign N126 = N123 | N125;
  assign N136 = N130 | N135;
  assign N149 = N143 | N148;
  assign N155 = N152 | N154;
  assign N156 = ~op_i[30];
  assign N164 = N161 | N163;
  assign N178 = N173 | N177;
  assign N179 = ~op_i[31];
  assign N180 = ~op_i[29];
  assign N181 = ~op_i[28];
  assign N182 = ~op_i[27];
  assign N183 = ~op_i[26];
  assign N184 = ~op_i[25];
  assign N214 = ~N213;
  assign N215 = N102 | N97;
  assign N216 = N108 | N215;
  assign N217 = N114 | N216;
  assign N218 = N120 | N217;
  assign N219 = N126 | N218;
  assign N220 = N136 | N219;
  assign N221 = N149 | N220;
  assign N222 = N155 | N221;
  assign N223 = N164 | N222;
  assign N224 = N178 | N223;
  assign N225 = N199 | N224;
  assign N226 = N207 | N225;
  assign N227 = N214 | N226;
  assign N228 = ~N227;
  assign N293 = ~carry;
  assign N294 = ~op_i[3];
  assign N300 = ~N299;
  assign N301 = ~op_i[13];
  assign N302 = ~op_i[12];
  assign N312 = ~op_i[14];
  assign N314 = ~rs1_eq_rs2;
  assign N315 = ~rs1_lt_rs2_signed;
  assign N316 = ~rs1_lt_rs2_unsigned;

endmodule



module bsg_dff_reset_en_width_p22_reset_val_p0_harden_p0
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [21:0] data_i;
  output [21:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [21:0] data_o;
  wire N0,N1,N2;
  reg data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = en_i;
  assign N1 = ~en_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_en_bypass_width_p22
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [21:0] data_i;
  output [21:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [21:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_reset_en_width_p22_reset_val_p0_harden_p0
  dff
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(en_i),
    .data_i(data_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_dff_en_width_p1
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input en_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_one_hot_width_p33_els_p3
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [98:0] data_i;
  input [2:0] sel_one_hot_i;
  output [32:0] data_o;
  wire [32:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32;
  wire [98:0] data_masked;
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[1];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[1];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[1];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[1];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[2];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[2];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[2];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[2];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[2];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[2];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[2];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[2];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[2];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[2];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[2];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[2];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[2];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[2];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[2];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[2];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[2];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[2];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[2];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[2];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[2];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[2];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[2];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[2];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[2];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[2];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[2];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[2];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[2];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[2];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[2];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[2];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[2];
  assign data_o[0] = N0 | data_masked[0];
  assign N0 = data_masked[66] | data_masked[33];
  assign data_o[1] = N1 | data_masked[1];
  assign N1 = data_masked[67] | data_masked[34];
  assign data_o[2] = N2 | data_masked[2];
  assign N2 = data_masked[68] | data_masked[35];
  assign data_o[3] = N3 | data_masked[3];
  assign N3 = data_masked[69] | data_masked[36];
  assign data_o[4] = N4 | data_masked[4];
  assign N4 = data_masked[70] | data_masked[37];
  assign data_o[5] = N5 | data_masked[5];
  assign N5 = data_masked[71] | data_masked[38];
  assign data_o[6] = N6 | data_masked[6];
  assign N6 = data_masked[72] | data_masked[39];
  assign data_o[7] = N7 | data_masked[7];
  assign N7 = data_masked[73] | data_masked[40];
  assign data_o[8] = N8 | data_masked[8];
  assign N8 = data_masked[74] | data_masked[41];
  assign data_o[9] = N9 | data_masked[9];
  assign N9 = data_masked[75] | data_masked[42];
  assign data_o[10] = N10 | data_masked[10];
  assign N10 = data_masked[76] | data_masked[43];
  assign data_o[11] = N11 | data_masked[11];
  assign N11 = data_masked[77] | data_masked[44];
  assign data_o[12] = N12 | data_masked[12];
  assign N12 = data_masked[78] | data_masked[45];
  assign data_o[13] = N13 | data_masked[13];
  assign N13 = data_masked[79] | data_masked[46];
  assign data_o[14] = N14 | data_masked[14];
  assign N14 = data_masked[80] | data_masked[47];
  assign data_o[15] = N15 | data_masked[15];
  assign N15 = data_masked[81] | data_masked[48];
  assign data_o[16] = N16 | data_masked[16];
  assign N16 = data_masked[82] | data_masked[49];
  assign data_o[17] = N17 | data_masked[17];
  assign N17 = data_masked[83] | data_masked[50];
  assign data_o[18] = N18 | data_masked[18];
  assign N18 = data_masked[84] | data_masked[51];
  assign data_o[19] = N19 | data_masked[19];
  assign N19 = data_masked[85] | data_masked[52];
  assign data_o[20] = N20 | data_masked[20];
  assign N20 = data_masked[86] | data_masked[53];
  assign data_o[21] = N21 | data_masked[21];
  assign N21 = data_masked[87] | data_masked[54];
  assign data_o[22] = N22 | data_masked[22];
  assign N22 = data_masked[88] | data_masked[55];
  assign data_o[23] = N23 | data_masked[23];
  assign N23 = data_masked[89] | data_masked[56];
  assign data_o[24] = N24 | data_masked[24];
  assign N24 = data_masked[90] | data_masked[57];
  assign data_o[25] = N25 | data_masked[25];
  assign N25 = data_masked[91] | data_masked[58];
  assign data_o[26] = N26 | data_masked[26];
  assign N26 = data_masked[92] | data_masked[59];
  assign data_o[27] = N27 | data_masked[27];
  assign N27 = data_masked[93] | data_masked[60];
  assign data_o[28] = N28 | data_masked[28];
  assign N28 = data_masked[94] | data_masked[61];
  assign data_o[29] = N29 | data_masked[29];
  assign N29 = data_masked[95] | data_masked[62];
  assign data_o[30] = N30 | data_masked[30];
  assign N30 = data_masked[96] | data_masked[63];
  assign data_o[31] = N31 | data_masked[31];
  assign N31 = data_masked[97] | data_masked[64];
  assign data_o[32] = N32 | data_masked[32];
  assign N32 = data_masked[98] | data_masked[65];

endmodule



module bsg_dff_en_width_p33
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [32:0] data_i;
  output [32:0] data_o;
  input clk_i;
  input en_i;
  wire [32:0] data_o;
  reg data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,
  data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,
  data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,
  data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_adder_cin_width_p33
(
  a_i,
  b_i,
  cin_i,
  o
);

  input [32:0] a_i;
  input [32:0] b_i;
  output [32:0] o;
  input cin_i;
  wire [32:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32;
  assign { N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } = a_i + b_i;
  assign o = { N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } + cin_i;

endmodule



module bsg_counter_clear_up_max_val_p32_init_val_p0_disable_overflow_warning_p1
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [5:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [5:0] count_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;
  reg count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,count_o_2_sv2v_reg,
  count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N12 = reset_i | clear_i;
  assign { N10, N9, N8, N7, N6, N5 } = count_o + up_i;
  assign N11 = (N0)? up_i : 
               (N1)? N5 : 1'b0;
  assign N0 = clear_i;
  assign N1 = N4;
  assign N2 = ~reset_i;
  assign N3 = N2;
  assign N4 = ~clear_i;

  always @(posedge clk_i) begin
    if(N12) begin
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_5_sv2v_reg <= N10;
      count_o_4_sv2v_reg <= N9;
      count_o_3_sv2v_reg <= N8;
      count_o_2_sv2v_reg <= N7;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_0_sv2v_reg <= N11;
    end 
  end


endmodule



module bsg_idiv_iterative_controller_width_p32
(
  clk_i,
  reset_i,
  v_i,
  ready_and_o,
  zero_divisor_i,
  signed_div_r_i,
  adder_result_is_neg_i,
  opA_is_neg_i,
  opC_is_neg_i,
  opA_sel_o,
  opA_ld_o,
  opA_inv_o,
  opA_clr_l_o,
  opB_sel_o,
  opB_ld_o,
  opB_inv_o,
  opB_clr_l_o,
  opC_sel_o,
  opC_ld_o,
  latch_signed_div_o,
  adder_cin_o,
  v_o,
  yumi_i
);

  output [2:0] opB_sel_o;
  output [2:0] opC_sel_o;
  input clk_i;
  input reset_i;
  input v_i;
  input zero_divisor_i;
  input signed_div_r_i;
  input adder_result_is_neg_i;
  input opA_is_neg_i;
  input opC_is_neg_i;
  input yumi_i;
  output ready_and_o;
  output opA_sel_o;
  output opA_ld_o;
  output opA_inv_o;
  output opA_clr_l_o;
  output opB_ld_o;
  output opB_inv_o;
  output opB_clr_l_o;
  output opC_ld_o;
  output latch_signed_div_o;
  output adder_cin_o;
  output v_o;
  wire [2:0] opB_sel_o,opC_sel_o;
  wire ready_and_o,opA_sel_o,opA_ld_o,opA_inv_o,opA_clr_l_o,opB_ld_o,opB_inv_o,
  opB_clr_l_o,opC_ld_o,latch_signed_div_o,adder_cin_o,v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,
  N10,N11,add_neg_last,neg_ld,N12,q_neg,N13,r_neg,calc_up_li,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N101,N102,N103,N104,N105,N106,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123;
  wire [5:0] state,calc_cnt;
  wire [3:0] next_state;
  reg add_neg_last_sv2v_reg,r_neg_sv2v_reg,q_neg_sv2v_reg,state_5_sv2v_reg,
  state_4_sv2v_reg,state_3_sv2v_reg,state_2_sv2v_reg,state_1_sv2v_reg,state_0_sv2v_reg;
  assign add_neg_last = add_neg_last_sv2v_reg;
  assign r_neg = r_neg_sv2v_reg;
  assign q_neg = q_neg_sv2v_reg;
  assign state[5] = state_5_sv2v_reg;
  assign state[4] = state_4_sv2v_reg;
  assign state[3] = state_3_sv2v_reg;
  assign state[2] = state_2_sv2v_reg;
  assign state[1] = state_1_sv2v_reg;
  assign state[0] = state_0_sv2v_reg;

  bsg_counter_clear_up_max_val_p32_init_val_p0_disable_overflow_warning_p1
  calc_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(N121),
    .up_i(calc_up_li),
    .count_o(calc_cnt)
  );

  assign N17 = N15 & N16;
  assign N20 = N101 & N108;
  assign N21 = N18 & N19;
  assign N22 = N20 & N21;
  assign N23 = state[3] | state[2];
  assign N24 = state[1] | N19;
  assign N25 = N23 | N24;
  assign N27 = state[3] | state[2];
  assign N28 = N18 | state[0];
  assign N29 = N27 | N28;
  assign N31 = state[3] | state[2];
  assign N32 = N18 | N19;
  assign N33 = N31 | N32;
  assign N35 = state[3] | N108;
  assign N36 = state[1] | state[0];
  assign N37 = N35 | N36;
  assign N39 = state[3] | N108;
  assign N40 = state[1] | N19;
  assign N41 = N39 | N40;
  assign N43 = state[3] | N108;
  assign N44 = N18 | state[0];
  assign N45 = N43 | N44;
  assign N47 = state[3] | N108;
  assign N48 = N18 | N19;
  assign N49 = N47 | N48;
  assign N51 = N101 | state[2];
  assign N52 = state[1] | state[0];
  assign N53 = N51 | N52;
  assign N95 = state[4] | state[5];
  assign N96 = state[3] | N95;
  assign N97 = state[2] | N96;
  assign N98 = state[1] | N97;
  assign N99 = state[0] | N98;
  assign ready_and_o = ~N99;
  assign N101 = ~state[3];
  assign N102 = state[4] | state[5];
  assign N103 = N101 | N102;
  assign N104 = state[2] | N103;
  assign N105 = state[1] | N104;
  assign N106 = state[0] | N105;
  assign v_o = ~N106;
  assign N108 = ~state[2];
  assign N109 = state[4] | state[5];
  assign N110 = state[3] | N109;
  assign N111 = N108 | N110;
  assign N112 = state[1] | N111;
  assign N113 = state[0] | N112;
  assign N114 = ~N113;
  assign N115 = ~calc_cnt[5];
  assign N116 = calc_cnt[4] | N115;
  assign N117 = calc_cnt[3] | N116;
  assign N118 = calc_cnt[2] | N117;
  assign N119 = calc_cnt[1] | N118;
  assign N120 = calc_cnt[0] | N119;
  assign N121 = ~N120;
  assign N55 = ~N13;
  assign { N61, N60 } = (N0)? { N59, adder_result_is_neg_i } : 
                        (N1)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = N58;
  assign N1 = N57;
  assign N63 = ~N62;
  assign { N77, N76, N75, N74 } = (N2)? { 1'b0, 1'b0, 1'b0, v_i } : 
                                  (N3)? { 1'b0, 1'b0, 1'b1, N55 } : 
                                  (N4)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                  (N5)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                  (N6)? { 1'b0, 1'b1, N61, N60 } : 
                                  (N7)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                  (N8)? { N62, N63, N63, N63 } : 
                                  (N9)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                  (N10)? { N64, 1'b0, 1'b0, 1'b0 } : 
                                  (N73)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N22;
  assign N3 = N26;
  assign N4 = N30;
  assign N5 = N34;
  assign N6 = N38;
  assign N7 = N42;
  assign N8 = N46;
  assign N9 = N50;
  assign N10 = N54;
  assign N78 = (N2)? v_i : 
               (N3)? N56 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b1 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N73)? 1'b0 : 1'b0;
  assign N79 = (N2)? 1'b1 : 
               (N3)? 1'b0 : 
               (N4)? 1'b1 : 
               (N5)? 1'b1 : 
               (N6)? 1'b1 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b1 : 
               (N10)? 1'b0 : 
               (N73)? 1'b1 : 1'b0;
  assign N80 = (N2)? v_i : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N73)? 1'b0 : 1'b0;
  assign N81 = (N2)? 1'b1 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N73)? 1'b0 : 1'b0;
  assign { N83, N82 } = (N2)? { 1'b0, 1'b0 } : 
                        (N3)? { 1'b0, 1'b1 } : 
                        (N4)? { 1'b1, 1'b0 } : 
                        (N5)? { 1'b0, 1'b1 } : 
                        (N6)? { 1'b0, 1'b1 } : 
                        (N7)? { 1'b0, 1'b1 } : 
                        (N8)? { 1'b0, 1'b1 } : 
                        (N9)? { 1'b1, 1'b0 } : 
                        (N10)? { 1'b0, 1'b1 } : 
                        (N73)? { 1'b0, 1'b1 } : 1'b0;
  assign N84 = (N2)? N14 : 
               (N3)? 1'b1 : 
               (N4)? N14 : 
               (N5)? N14 : 
               (N6)? N14 : 
               (N7)? 1'b0 : 
               (N8)? N14 : 
               (N9)? N14 : 
               (N10)? N14 : 
               (N73)? N14 : 1'b0;
  assign N85 = (N2)? 1'b1 : 
               (N3)? 1'b0 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N6)? 1'b1 : 
               (N7)? 1'b1 : 
               (N8)? 1'b1 : 
               (N9)? 1'b1 : 
               (N10)? 1'b1 : 
               (N73)? 1'b1 : 1'b0;
  assign { N88, N87, N86 } = (N2)? { 1'b0, 1'b0, 1'b1 } : 
                             (N3)? { 1'b1, 1'b0, 1'b0 } : 
                             (N4)? { 1'b0, 1'b0, 1'b1 } : 
                             (N5)? { 1'b0, 1'b0, 1'b1 } : 
                             (N6)? { 1'b0, N58, N57 } : 
                             (N7)? { 1'b0, 1'b1, 1'b0 } : 
                             (N8)? { 1'b1, 1'b0, 1'b0 } : 
                             (N9)? { 1'b0, 1'b0, 1'b1 } : 
                             (N10)? { 1'b0, 1'b0, 1'b1 } : 
                             (N73)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign N89 = (N2)? 1'b0 : 
               (N3)? 1'b1 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N73)? 1'b0 : 1'b0;
  assign N90 = (N2)? N14 : 
               (N3)? 1'b1 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N6)? N14 : 
               (N7)? 1'b0 : 
               (N8)? r_neg : 
               (N9)? 1'b1 : 
               (N10)? N14 : 
               (N73)? N14 : 1'b0;
  assign N91 = (N2)? 1'b1 : 
               (N3)? 1'b1 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N6)? 1'b1 : 
               (N7)? 1'b1 : 
               (N8)? 1'b0 : 
               (N9)? 1'b0 : 
               (N10)? 1'b1 : 
               (N73)? 1'b1 : 1'b0;
  assign N92 = (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N8)? r_neg : 
               (N9)? 1'b1 : 
               (N10)? 1'b0 : 
               (N73)? 1'b0 : 1'b0;
  assign N93 = (N2)? 1'b1 : 
               (N3)? 1'b1 : 
               (N4)? 1'b0 : 
               (N5)? 1'b1 : 
               (N6)? 1'b1 : 
               (N7)? 1'b1 : 
               (N8)? 1'b1 : 
               (N9)? 1'b0 : 
               (N10)? 1'b0 : 
               (N73)? 1'b1 : 1'b0;
  assign opB_inv_o = (N11)? N92 : 
                     (N94)? 1'b0 : 1'b0;
  assign N11 = N17;
  assign opB_ld_o = (N11)? N93 : 
                    (N94)? 1'b1 : 1'b0;
  assign next_state = (N11)? { N77, N76, N75, N74 } : 
                      (N94)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign opA_ld_o = (N11)? N78 : 
                    (N94)? 1'b0 : 1'b0;
  assign opC_ld_o = (N11)? N79 : 
                    (N94)? 1'b1 : 1'b0;
  assign latch_signed_div_o = (N11)? N80 : 
                              (N94)? 1'b0 : 1'b0;
  assign opA_sel_o = (N11)? N81 : 
                     (N94)? 1'b0 : 1'b0;
  assign opC_sel_o = (N11)? { N22, N83, N82 } : 
                     (N94)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign opA_inv_o = (N11)? N84 : 
                     (N94)? N14 : 1'b0;
  assign opB_clr_l_o = (N11)? N85 : 
                       (N94)? 1'b1 : 1'b0;
  assign opB_sel_o = (N11)? { N88, N87, N86 } : 
                     (N94)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign neg_ld = (N11)? N89 : 
                  (N94)? 1'b0 : 1'b0;
  assign adder_cin_o = (N11)? N90 : 
                       (N94)? N14 : 1'b0;
  assign opA_clr_l_o = (N11)? N91 : 
                       (N94)? 1'b1 : 1'b0;
  assign N12 = N122 & signed_div_r_i;
  assign N122 = opA_is_neg_i ^ opC_is_neg_i;
  assign N13 = opC_is_neg_i & signed_div_r_i;
  assign calc_up_li = N114 & N115;
  assign N14 = ~add_neg_last;
  assign N15 = ~state[5];
  assign N16 = ~state[4];
  assign N18 = ~state[1];
  assign N19 = ~state[0];
  assign N26 = ~N25;
  assign N30 = ~N29;
  assign N34 = ~N33;
  assign N38 = ~N37;
  assign N42 = ~N41;
  assign N46 = ~N45;
  assign N50 = ~N49;
  assign N54 = ~N53;
  assign N56 = opA_is_neg_i & signed_div_r_i;
  assign N57 = ~N121;
  assign N58 = N121;
  assign N59 = ~adder_result_is_neg_i;
  assign N62 = zero_divisor_i | N123;
  assign N123 = ~q_neg;
  assign N64 = ~yumi_i;
  assign N65 = N26 | N22;
  assign N66 = N30 | N65;
  assign N67 = N34 | N66;
  assign N68 = N38 | N67;
  assign N69 = N42 | N68;
  assign N70 = N46 | N69;
  assign N71 = N50 | N70;
  assign N72 = N54 | N71;
  assign N73 = ~N72;
  assign N94 = ~N17;

  always @(posedge clk_i) begin
    if(1'b1) begin
      add_neg_last_sv2v_reg <= adder_result_is_neg_i;
    end 
    if(neg_ld) begin
      r_neg_sv2v_reg <= N13;
      q_neg_sv2v_reg <= N12;
    end 
    if(reset_i) begin
      state_5_sv2v_reg <= 1'b0;
      state_4_sv2v_reg <= 1'b0;
      state_3_sv2v_reg <= 1'b0;
      state_2_sv2v_reg <= 1'b0;
      state_1_sv2v_reg <= 1'b0;
      state_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      state_5_sv2v_reg <= 1'b0;
      state_4_sv2v_reg <= 1'b0;
      state_3_sv2v_reg <= next_state[3];
      state_2_sv2v_reg <= next_state[2];
      state_1_sv2v_reg <= next_state[1];
      state_0_sv2v_reg <= next_state[0];
    end 
  end


endmodule



module bsg_idiv_iterative
(
  clk_i,
  reset_i,
  v_i,
  ready_and_o,
  dividend_i,
  divisor_i,
  signed_div_i,
  v_o,
  quotient_o,
  remainder_o,
  yumi_i
);

  input [31:0] dividend_i;
  input [31:0] divisor_i;
  output [31:0] quotient_o;
  output [31:0] remainder_o;
  input clk_i;
  input reset_i;
  input v_i;
  input signed_div_i;
  input yumi_i;
  output ready_and_o;
  output v_o;
  wire [31:0] quotient_o,remainder_o;
  wire ready_and_o,v_o,divisor_msb,dividend_msb,signed_div_r,latch_signed_div_lo,
  zero_divisor_li,opA_sel_lo,_2_net__0_,opA_ld_lo,opB_ld_lo,opC_ld_lo,opA_inv_lo,
  opA_clr_lo,opB_inv_lo,opB_clr_lo,adder_cin_lo,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97;
  wire [32:32] opA_r,opC_r;
  wire [32:0] opA_mux,add_out,opB_mux,opC_mux,opB_r,add_in0,add_in1;
  wire [2:0] opB_sel_lo,opC_sel_lo;

  bsg_dff_en_width_p1
  req_reg
  (
    .clk_i(clk_i),
    .data_i(signed_div_i),
    .en_i(latch_signed_div_lo),
    .data_o(signed_div_r)
  );


  bsg_mux_width_p33_els_p2
  muxA
  (
    .data_i({ divisor_msb, divisor_i, add_out }),
    .sel_i(opA_sel_lo),
    .data_o(opA_mux)
  );


  bsg_mux_one_hot_width_p33_els_p3
  muxB
  (
    .data_i({ opC_r[32:32], quotient_o, add_out, add_out[31:0], opC_r[32:32] }),
    .sel_one_hot_i(opB_sel_lo),
    .data_o(opB_mux)
  );


  bsg_mux_one_hot_width_p33_els_p3
  muxC
  (
    .data_i({ dividend_msb, dividend_i, add_out, quotient_o, _2_net__0_ }),
    .sel_one_hot_i(opC_sel_lo),
    .data_o(opC_mux)
  );


  bsg_dff_en_width_p33
  opA_reg
  (
    .clk_i(clk_i),
    .data_i(opA_mux),
    .en_i(opA_ld_lo),
    .data_o({ opA_r[32:32], remainder_o })
  );


  bsg_dff_en_width_p33
  opB_reg
  (
    .clk_i(clk_i),
    .data_i(opB_mux),
    .en_i(opB_ld_lo),
    .data_o(opB_r)
  );


  bsg_dff_en_width_p33
  opC_reg
  (
    .clk_i(clk_i),
    .data_i(opC_mux),
    .en_i(opC_ld_lo),
    .data_o({ opC_r[32:32], quotient_o })
  );


  bsg_adder_cin_width_p33
  adder
  (
    .a_i(add_in0),
    .b_i(add_in1),
    .cin_i(adder_cin_lo),
    .o(add_out)
  );


  bsg_idiv_iterative_controller_width_p32
  control
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_and_o(ready_and_o),
    .zero_divisor_i(zero_divisor_li),
    .signed_div_r_i(signed_div_r),
    .adder_result_is_neg_i(add_out[32]),
    .opA_is_neg_i(opA_r[32]),
    .opC_is_neg_i(opC_r[32]),
    .opA_sel_o(opA_sel_lo),
    .opA_ld_o(opA_ld_lo),
    .opA_inv_o(opA_inv_lo),
    .opA_clr_l_o(opA_clr_lo),
    .opB_sel_o(opB_sel_lo),
    .opB_ld_o(opB_ld_lo),
    .opB_inv_o(opB_inv_lo),
    .opB_clr_l_o(opB_clr_lo),
    .opC_sel_o(opC_sel_lo),
    .opC_ld_o(opC_ld_lo),
    .latch_signed_div_o(latch_signed_div_lo),
    .adder_cin_o(adder_cin_lo),
    .v_o(v_o),
    .yumi_i(yumi_i)
  );

  assign divisor_msb = signed_div_i & divisor_i[31];
  assign dividend_msb = signed_div_i & dividend_i[31];
  assign zero_divisor_li = ~N31;
  assign N31 = N30 | remainder_o[0];
  assign N30 = N29 | remainder_o[1];
  assign N29 = N28 | remainder_o[2];
  assign N28 = N27 | remainder_o[3];
  assign N27 = N26 | remainder_o[4];
  assign N26 = N25 | remainder_o[5];
  assign N25 = N24 | remainder_o[6];
  assign N24 = N23 | remainder_o[7];
  assign N23 = N22 | remainder_o[8];
  assign N22 = N21 | remainder_o[9];
  assign N21 = N20 | remainder_o[10];
  assign N20 = N19 | remainder_o[11];
  assign N19 = N18 | remainder_o[12];
  assign N18 = N17 | remainder_o[13];
  assign N17 = N16 | remainder_o[14];
  assign N16 = N15 | remainder_o[15];
  assign N15 = N14 | remainder_o[16];
  assign N14 = N13 | remainder_o[17];
  assign N13 = N12 | remainder_o[18];
  assign N12 = N11 | remainder_o[19];
  assign N11 = N10 | remainder_o[20];
  assign N10 = N9 | remainder_o[21];
  assign N9 = N8 | remainder_o[22];
  assign N8 = N7 | remainder_o[23];
  assign N7 = N6 | remainder_o[24];
  assign N6 = N5 | remainder_o[25];
  assign N5 = N4 | remainder_o[26];
  assign N4 = N3 | remainder_o[27];
  assign N3 = N2 | remainder_o[28];
  assign N2 = N1 | remainder_o[29];
  assign N1 = N0 | remainder_o[30];
  assign N0 = opA_r[32] | remainder_o[31];
  assign _2_net__0_ = ~add_out[32];
  assign add_in0[32] = N32 & opA_clr_lo;
  assign N32 = opA_r[32] ^ opA_inv_lo;
  assign add_in0[31] = N33 & opA_clr_lo;
  assign N33 = remainder_o[31] ^ opA_inv_lo;
  assign add_in0[30] = N34 & opA_clr_lo;
  assign N34 = remainder_o[30] ^ opA_inv_lo;
  assign add_in0[29] = N35 & opA_clr_lo;
  assign N35 = remainder_o[29] ^ opA_inv_lo;
  assign add_in0[28] = N36 & opA_clr_lo;
  assign N36 = remainder_o[28] ^ opA_inv_lo;
  assign add_in0[27] = N37 & opA_clr_lo;
  assign N37 = remainder_o[27] ^ opA_inv_lo;
  assign add_in0[26] = N38 & opA_clr_lo;
  assign N38 = remainder_o[26] ^ opA_inv_lo;
  assign add_in0[25] = N39 & opA_clr_lo;
  assign N39 = remainder_o[25] ^ opA_inv_lo;
  assign add_in0[24] = N40 & opA_clr_lo;
  assign N40 = remainder_o[24] ^ opA_inv_lo;
  assign add_in0[23] = N41 & opA_clr_lo;
  assign N41 = remainder_o[23] ^ opA_inv_lo;
  assign add_in0[22] = N42 & opA_clr_lo;
  assign N42 = remainder_o[22] ^ opA_inv_lo;
  assign add_in0[21] = N43 & opA_clr_lo;
  assign N43 = remainder_o[21] ^ opA_inv_lo;
  assign add_in0[20] = N44 & opA_clr_lo;
  assign N44 = remainder_o[20] ^ opA_inv_lo;
  assign add_in0[19] = N45 & opA_clr_lo;
  assign N45 = remainder_o[19] ^ opA_inv_lo;
  assign add_in0[18] = N46 & opA_clr_lo;
  assign N46 = remainder_o[18] ^ opA_inv_lo;
  assign add_in0[17] = N47 & opA_clr_lo;
  assign N47 = remainder_o[17] ^ opA_inv_lo;
  assign add_in0[16] = N48 & opA_clr_lo;
  assign N48 = remainder_o[16] ^ opA_inv_lo;
  assign add_in0[15] = N49 & opA_clr_lo;
  assign N49 = remainder_o[15] ^ opA_inv_lo;
  assign add_in0[14] = N50 & opA_clr_lo;
  assign N50 = remainder_o[14] ^ opA_inv_lo;
  assign add_in0[13] = N51 & opA_clr_lo;
  assign N51 = remainder_o[13] ^ opA_inv_lo;
  assign add_in0[12] = N52 & opA_clr_lo;
  assign N52 = remainder_o[12] ^ opA_inv_lo;
  assign add_in0[11] = N53 & opA_clr_lo;
  assign N53 = remainder_o[11] ^ opA_inv_lo;
  assign add_in0[10] = N54 & opA_clr_lo;
  assign N54 = remainder_o[10] ^ opA_inv_lo;
  assign add_in0[9] = N55 & opA_clr_lo;
  assign N55 = remainder_o[9] ^ opA_inv_lo;
  assign add_in0[8] = N56 & opA_clr_lo;
  assign N56 = remainder_o[8] ^ opA_inv_lo;
  assign add_in0[7] = N57 & opA_clr_lo;
  assign N57 = remainder_o[7] ^ opA_inv_lo;
  assign add_in0[6] = N58 & opA_clr_lo;
  assign N58 = remainder_o[6] ^ opA_inv_lo;
  assign add_in0[5] = N59 & opA_clr_lo;
  assign N59 = remainder_o[5] ^ opA_inv_lo;
  assign add_in0[4] = N60 & opA_clr_lo;
  assign N60 = remainder_o[4] ^ opA_inv_lo;
  assign add_in0[3] = N61 & opA_clr_lo;
  assign N61 = remainder_o[3] ^ opA_inv_lo;
  assign add_in0[2] = N62 & opA_clr_lo;
  assign N62 = remainder_o[2] ^ opA_inv_lo;
  assign add_in0[1] = N63 & opA_clr_lo;
  assign N63 = remainder_o[1] ^ opA_inv_lo;
  assign add_in0[0] = N64 & opA_clr_lo;
  assign N64 = remainder_o[0] ^ opA_inv_lo;
  assign add_in1[32] = N65 & opB_clr_lo;
  assign N65 = opB_r[32] ^ opB_inv_lo;
  assign add_in1[31] = N66 & opB_clr_lo;
  assign N66 = opB_r[31] ^ opB_inv_lo;
  assign add_in1[30] = N67 & opB_clr_lo;
  assign N67 = opB_r[30] ^ opB_inv_lo;
  assign add_in1[29] = N68 & opB_clr_lo;
  assign N68 = opB_r[29] ^ opB_inv_lo;
  assign add_in1[28] = N69 & opB_clr_lo;
  assign N69 = opB_r[28] ^ opB_inv_lo;
  assign add_in1[27] = N70 & opB_clr_lo;
  assign N70 = opB_r[27] ^ opB_inv_lo;
  assign add_in1[26] = N71 & opB_clr_lo;
  assign N71 = opB_r[26] ^ opB_inv_lo;
  assign add_in1[25] = N72 & opB_clr_lo;
  assign N72 = opB_r[25] ^ opB_inv_lo;
  assign add_in1[24] = N73 & opB_clr_lo;
  assign N73 = opB_r[24] ^ opB_inv_lo;
  assign add_in1[23] = N74 & opB_clr_lo;
  assign N74 = opB_r[23] ^ opB_inv_lo;
  assign add_in1[22] = N75 & opB_clr_lo;
  assign N75 = opB_r[22] ^ opB_inv_lo;
  assign add_in1[21] = N76 & opB_clr_lo;
  assign N76 = opB_r[21] ^ opB_inv_lo;
  assign add_in1[20] = N77 & opB_clr_lo;
  assign N77 = opB_r[20] ^ opB_inv_lo;
  assign add_in1[19] = N78 & opB_clr_lo;
  assign N78 = opB_r[19] ^ opB_inv_lo;
  assign add_in1[18] = N79 & opB_clr_lo;
  assign N79 = opB_r[18] ^ opB_inv_lo;
  assign add_in1[17] = N80 & opB_clr_lo;
  assign N80 = opB_r[17] ^ opB_inv_lo;
  assign add_in1[16] = N81 & opB_clr_lo;
  assign N81 = opB_r[16] ^ opB_inv_lo;
  assign add_in1[15] = N82 & opB_clr_lo;
  assign N82 = opB_r[15] ^ opB_inv_lo;
  assign add_in1[14] = N83 & opB_clr_lo;
  assign N83 = opB_r[14] ^ opB_inv_lo;
  assign add_in1[13] = N84 & opB_clr_lo;
  assign N84 = opB_r[13] ^ opB_inv_lo;
  assign add_in1[12] = N85 & opB_clr_lo;
  assign N85 = opB_r[12] ^ opB_inv_lo;
  assign add_in1[11] = N86 & opB_clr_lo;
  assign N86 = opB_r[11] ^ opB_inv_lo;
  assign add_in1[10] = N87 & opB_clr_lo;
  assign N87 = opB_r[10] ^ opB_inv_lo;
  assign add_in1[9] = N88 & opB_clr_lo;
  assign N88 = opB_r[9] ^ opB_inv_lo;
  assign add_in1[8] = N89 & opB_clr_lo;
  assign N89 = opB_r[8] ^ opB_inv_lo;
  assign add_in1[7] = N90 & opB_clr_lo;
  assign N90 = opB_r[7] ^ opB_inv_lo;
  assign add_in1[6] = N91 & opB_clr_lo;
  assign N91 = opB_r[6] ^ opB_inv_lo;
  assign add_in1[5] = N92 & opB_clr_lo;
  assign N92 = opB_r[5] ^ opB_inv_lo;
  assign add_in1[4] = N93 & opB_clr_lo;
  assign N93 = opB_r[4] ^ opB_inv_lo;
  assign add_in1[3] = N94 & opB_clr_lo;
  assign N94 = opB_r[3] ^ opB_inv_lo;
  assign add_in1[2] = N95 & opB_clr_lo;
  assign N95 = opB_r[2] ^ opB_inv_lo;
  assign add_in1[1] = N96 & opB_clr_lo;
  assign N96 = opB_r[1] ^ opB_inv_lo;
  assign add_in1[0] = N97 & opB_clr_lo;
  assign N97 = opB_r[0] ^ opB_inv_lo;

endmodule



module idiv
(
  clk_i,
  reset_i,
  v_i,
  rs1_i,
  rs2_i,
  rd_i,
  op_i,
  ready_o,
  v_o,
  rd_o,
  result_o,
  yumi_i
);

  input [31:0] rs1_i;
  input [31:0] rs2_i;
  input [4:0] rd_i;
  input [1:0] op_i;
  output [4:0] rd_o;
  output [31:0] result_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [4:0] rd_o;
  wire [31:0] result_o,quotient_lo,remainder_lo;
  wire ready_o,v_o,N0,N1,N3,signed_div_li,N4,rem_r,N5,N6,N7,N2,N8,N9,N10,N11,N12,N13;
  reg rem_r_sv2v_reg,rd_o_4_sv2v_reg,rd_o_3_sv2v_reg,rd_o_2_sv2v_reg,rd_o_1_sv2v_reg,
  rd_o_0_sv2v_reg;
  assign rem_r = rem_r_sv2v_reg;
  assign rd_o[4] = rd_o_4_sv2v_reg;
  assign rd_o[3] = rd_o_3_sv2v_reg;
  assign rd_o[2] = rd_o_2_sv2v_reg;
  assign rd_o[1] = rd_o_1_sv2v_reg;
  assign rd_o[0] = rd_o_0_sv2v_reg;

  bsg_idiv_iterative
  idiv0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_and_o(ready_o),
    .dividend_i(rs1_i),
    .divisor_i(rs2_i),
    .signed_div_i(signed_div_li),
    .v_o(v_o),
    .quotient_o(quotient_lo),
    .remainder_o(remainder_lo),
    .yumi_i(yumi_i)
  );

  assign N8 = op_i[0] | op_i[1];
  assign N9 = ~N8;
  assign N10 = ~op_i[1];
  assign N11 = op_i[0] | N10;
  assign N12 = ~N11;
  assign N13 = op_i[0] & op_i[1];
  assign N6 = (N0)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = N4;
  assign result_o = (N1)? remainder_lo : 
                    (N3)? quotient_lo : 1'b0;
  assign N1 = rem_r;
  assign N3 = N7;
  assign signed_div_li = N12 | N9;
  assign N4 = v_i & ready_o;
  assign N5 = N12 | N13;
  assign N7 = ~rem_r;
  assign N2 = ~N4;

  always @(posedge clk_i) begin
    if(reset_i) begin
      rem_r_sv2v_reg <= 1'b0;
      rd_o_4_sv2v_reg <= 1'b0;
      rd_o_3_sv2v_reg <= 1'b0;
      rd_o_2_sv2v_reg <= 1'b0;
      rd_o_1_sv2v_reg <= 1'b0;
      rd_o_0_sv2v_reg <= 1'b0;
    end else if(N6) begin
      rem_r_sv2v_reg <= N5;
      rd_o_4_sv2v_reg <= rd_i[4];
      rd_o_3_sv2v_reg <= rd_i[3];
      rd_o_2_sv2v_reg <= rd_i[2];
      rd_o_1_sv2v_reg <= rd_i[1];
      rd_o_0_sv2v_reg <= rd_i[0];
    end 
  end


endmodule



module lsu_data_width_p32_pc_width_p22_dmem_size_p1024
(
  clk_i,
  reset_i,
  exe_decode_i,
  exe_rs1_i,
  exe_rs2_i,
  exe_rd_i,
  mem_offset_i,
  pc_plus4_i,
  icache_miss_i,
  remote_req_o,
  remote_req_v_o,
  dmem_v_o,
  dmem_w_o,
  dmem_addr_o,
  dmem_data_o,
  dmem_mask_o,
  reserve_o,
  mem_addr_sent_o
);

  input [30:0] exe_decode_i;
  input [31:0] exe_rs1_i;
  input [31:0] exe_rs2_i;
  input [4:0] exe_rd_i;
  input [31:0] mem_offset_i;
  input [31:0] pc_plus4_i;
  output [83:0] remote_req_o;
  output [9:0] dmem_addr_o;
  output [31:0] dmem_data_o;
  output [3:0] dmem_mask_o;
  output [31:0] mem_addr_sent_o;
  input clk_i;
  input reset_i;
  input icache_miss_i;
  output remote_req_v_o;
  output dmem_v_o;
  output dmem_w_o;
  output reserve_o;
  wire [83:0] remote_req_o;
  wire [9:0] dmem_addr_o;
  wire [31:0] dmem_data_o,mem_addr_sent_o;
  wire [3:0] dmem_mask_o;
  wire remote_req_v_o,dmem_v_o,dmem_w_o,reserve_o,N0,N1,N2,
  remote_req_o_write_not_read_,remote_req_o_is_amo_op_,remote_req_o_amo_type__1_,remote_req_o_amo_type__0_,
  remote_req_o_reg_id__4_,remote_req_o_reg_id__3_,remote_req_o_reg_id__2_,
  remote_req_o_reg_id__1_,remote_req_o_reg_id__0_,mem_addr_1,mem_addr_0,N3,N4,N5,N6,N7,N8,N9,
  N10,is_local_dmem_addr,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58;
  wire [31:12] mem_addr;
  wire [30:0] miss_addr;
  assign remote_req_o_write_not_read_ = exe_decode_i[26];
  assign dmem_w_o = remote_req_o_write_not_read_;
  assign remote_req_o[83] = remote_req_o_write_not_read_;
  assign remote_req_o_is_amo_op_ = exe_decode_i[12];
  assign remote_req_o[82] = remote_req_o_is_amo_op_;
  assign remote_req_o_amo_type__1_ = exe_decode_i[9];
  assign remote_req_o[81] = remote_req_o_amo_type__1_;
  assign remote_req_o_amo_type__0_ = exe_decode_i[8];
  assign remote_req_o[80] = remote_req_o_amo_type__0_;
  assign remote_req_o_reg_id__4_ = exe_rd_i[4];
  assign remote_req_o[68] = remote_req_o_reg_id__4_;
  assign remote_req_o_reg_id__3_ = exe_rd_i[3];
  assign remote_req_o[67] = remote_req_o_reg_id__3_;
  assign remote_req_o_reg_id__2_ = exe_rd_i[2];
  assign remote_req_o[66] = remote_req_o_reg_id__2_;
  assign remote_req_o_reg_id__1_ = exe_rd_i[1];
  assign remote_req_o[65] = remote_req_o_reg_id__1_;
  assign remote_req_o_reg_id__0_ = exe_rd_i[0];
  assign remote_req_o[64] = remote_req_o_reg_id__0_;
  assign remote_req_o[63] = dmem_data_o[31];
  assign remote_req_o[62] = dmem_data_o[30];
  assign remote_req_o[61] = dmem_data_o[29];
  assign remote_req_o[60] = dmem_data_o[28];
  assign remote_req_o[59] = dmem_data_o[27];
  assign remote_req_o[58] = dmem_data_o[26];
  assign remote_req_o[57] = dmem_data_o[25];
  assign remote_req_o[56] = dmem_data_o[24];
  assign remote_req_o[55] = dmem_data_o[23];
  assign remote_req_o[54] = dmem_data_o[22];
  assign remote_req_o[53] = dmem_data_o[21];
  assign remote_req_o[52] = dmem_data_o[20];
  assign remote_req_o[51] = dmem_data_o[19];
  assign remote_req_o[50] = dmem_data_o[18];
  assign remote_req_o[49] = dmem_data_o[17];
  assign remote_req_o[48] = dmem_data_o[16];
  assign remote_req_o[47] = dmem_data_o[15];
  assign remote_req_o[46] = dmem_data_o[14];
  assign remote_req_o[45] = dmem_data_o[13];
  assign remote_req_o[44] = dmem_data_o[12];
  assign remote_req_o[43] = dmem_data_o[11];
  assign remote_req_o[42] = dmem_data_o[10];
  assign remote_req_o[41] = dmem_data_o[9];
  assign remote_req_o[40] = dmem_data_o[8];
  assign dmem_data_o[7] = exe_rs2_i[7];
  assign remote_req_o[39] = dmem_data_o[7];
  assign dmem_data_o[6] = exe_rs2_i[6];
  assign remote_req_o[38] = dmem_data_o[6];
  assign dmem_data_o[5] = exe_rs2_i[5];
  assign remote_req_o[37] = dmem_data_o[5];
  assign dmem_data_o[4] = exe_rs2_i[4];
  assign remote_req_o[36] = dmem_data_o[4];
  assign dmem_data_o[3] = exe_rs2_i[3];
  assign remote_req_o[35] = dmem_data_o[3];
  assign dmem_data_o[2] = exe_rs2_i[2];
  assign remote_req_o[34] = dmem_data_o[2];
  assign dmem_data_o[1] = exe_rs2_i[1];
  assign remote_req_o[33] = dmem_data_o[1];
  assign dmem_data_o[0] = exe_rs2_i[0];
  assign remote_req_o[32] = dmem_data_o[0];
  assign remote_req_o[79] = dmem_mask_o[3];
  assign remote_req_o[78] = dmem_mask_o[2];
  assign remote_req_o[77] = dmem_mask_o[1];
  assign remote_req_o[76] = dmem_mask_o[0];
  assign { mem_addr, dmem_addr_o, mem_addr_1, mem_addr_0 } = exe_rs1_i + mem_offset_i;
  assign miss_addr = pc_plus4_i[30:0] - { 1'b1, 1'b0, 1'b0 };
  assign dmem_data_o[31:8] = (N0)? { dmem_data_o[7:0], dmem_data_o[7:0], dmem_data_o[7:0] } : 
                             (N10)? { exe_rs2_i[15:8], dmem_data_o[7:0], exe_rs2_i[15:8] } : 
                             (N4)? exe_rs2_i[31:8] : 1'b0;
  assign N0 = exe_decode_i[25];
  assign dmem_mask_o = (N0)? { N5, N6, N7, N8 } : 
                       (N10)? { mem_addr_1, mem_addr_1, N13, N13 } : 
                       (N4)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign mem_addr_sent_o = (N1)? { 1'b1, miss_addr } : 
                           (N2)? { mem_addr, dmem_addr_o, mem_addr_1, mem_addr_0 } : 1'b0;
  assign N1 = remote_req_o[74];
  assign N2 = N11;
  assign { remote_req_o[75:75], remote_req_o[73:69] } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2)? { exe_decode_i[3:3], exe_decode_i[23:23], exe_decode_i[25:24], mem_addr_1, mem_addr_0 } : 1'b0;
  assign remote_req_o[31:0] = (N1)? { 1'b1, miss_addr } : 
                              (N2)? { mem_addr, dmem_addr_o, mem_addr_1, mem_addr_0 } : 1'b0;
  assign N3 = exe_decode_i[24] | exe_decode_i[25];
  assign N4 = ~N3;
  assign N5 = mem_addr_1 & mem_addr_0;
  assign N6 = mem_addr_1 & N12;
  assign N12 = ~mem_addr_0;
  assign N7 = N13 & mem_addr_0;
  assign N13 = ~mem_addr_1;
  assign N8 = N13 & N12;
  assign N9 = ~exe_decode_i[25];
  assign N10 = exe_decode_i[24] & N9;
  assign is_local_dmem_addr = N50 & N51;
  assign N50 = N48 & N49;
  assign N48 = N46 & N47;
  assign N46 = N44 & N45;
  assign N44 = N42 & N43;
  assign N42 = N40 & N41;
  assign N40 = N38 & N39;
  assign N38 = N36 & N37;
  assign N36 = N34 & N35;
  assign N34 = N32 & N33;
  assign N32 = N30 & N31;
  assign N30 = N28 & N29;
  assign N28 = N26 & N27;
  assign N26 = N24 & N25;
  assign N24 = N22 & N23;
  assign N22 = N20 & N21;
  assign N20 = N18 & N19;
  assign N18 = N16 & N17;
  assign N16 = N14 & N15;
  assign N14 = ~mem_addr[31];
  assign N15 = ~mem_addr[30];
  assign N17 = ~mem_addr[29];
  assign N19 = ~mem_addr[28];
  assign N21 = ~mem_addr[27];
  assign N23 = ~mem_addr[26];
  assign N25 = ~mem_addr[25];
  assign N27 = ~mem_addr[24];
  assign N29 = ~mem_addr[23];
  assign N31 = ~mem_addr[22];
  assign N33 = ~mem_addr[21];
  assign N35 = ~mem_addr[20];
  assign N37 = ~mem_addr[19];
  assign N39 = ~mem_addr[18];
  assign N41 = ~mem_addr[17];
  assign N43 = ~mem_addr[16];
  assign N45 = ~mem_addr[15];
  assign N47 = ~mem_addr[14];
  assign N49 = ~mem_addr[13];
  assign N51 = ~mem_addr[12];
  assign dmem_v_o = is_local_dmem_addr & N54;
  assign N54 = N53 | exe_decode_i[14];
  assign N53 = N52 | exe_decode_i[13];
  assign N52 = exe_decode_i[27] | remote_req_o_write_not_read_;
  assign N11 = ~icache_miss_i;
  assign remote_req_o[74] = icache_miss_i;
  assign remote_req_v_o = icache_miss_i | N58;
  assign N58 = N56 & N57;
  assign N56 = N55 | remote_req_o_is_amo_op_;
  assign N55 = exe_decode_i[27] | remote_req_o_write_not_read_;
  assign N57 = ~is_local_dmem_addr;
  assign reserve_o = exe_decode_i[13] & is_local_dmem_addr;

endmodule



module bsg_dff_en_width_p22_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [21:0] data_i;
  output [21:0] data_o;
  input clk_i;
  input en_i;
  wire [21:0] data_o;
  reg data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,
  data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,
  data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,
  data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,
  data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,
  data_o_0_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p22
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [21:0] data_i;
  output [21:0] data_o;
  input clk_i;
  input en_i;
  wire [21:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p22_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_dff_reset_width_p19
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [18:0] data_i;
  output [18:0] data_o;
  input clk_i;
  input reset_i;
  wire [18:0] data_o;
  reg data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p99
(
  clk_i,
  data_i,
  data_o
);

  input [98:0] data_i;
  output [98:0] data_o;
  input clk_i;
  wire [98:0] data_o;
  reg data_o_98_sv2v_reg,data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,
  data_o_94_sv2v_reg,data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,
  data_o_90_sv2v_reg,data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,
  data_o_86_sv2v_reg,data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,
  data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,
  data_o_77_sv2v_reg,data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,
  data_o_73_sv2v_reg,data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,
  data_o_69_sv2v_reg,data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,
  data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,
  data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,
  data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,
  data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,
  data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,
  data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,
  data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_98_sv2v_reg <= data_i[98];
      data_o_97_sv2v_reg <= data_i[97];
      data_o_96_sv2v_reg <= data_i[96];
      data_o_95_sv2v_reg <= data_i[95];
      data_o_94_sv2v_reg <= data_i[94];
      data_o_93_sv2v_reg <= data_i[93];
      data_o_92_sv2v_reg <= data_i[92];
      data_o_91_sv2v_reg <= data_i[91];
      data_o_90_sv2v_reg <= data_i[90];
      data_o_89_sv2v_reg <= data_i[89];
      data_o_88_sv2v_reg <= data_i[88];
      data_o_87_sv2v_reg <= data_i[87];
      data_o_86_sv2v_reg <= data_i[86];
      data_o_85_sv2v_reg <= data_i[85];
      data_o_84_sv2v_reg <= data_i[84];
      data_o_83_sv2v_reg <= data_i[83];
      data_o_82_sv2v_reg <= data_i[82];
      data_o_81_sv2v_reg <= data_i[81];
      data_o_80_sv2v_reg <= data_i[80];
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module isSigNaNRecFN_expWidth8_sigWidth24
(
  in,
  isSigNaN
);

  input [32:0] in;
  output isSigNaN;
  wire isSigNaN,N0,N1,N2;
  assign N0 = in[30] & in[31];
  assign N1 = in[29] & N0;
  assign isSigNaN = N1 & N2;
  assign N2 = ~in[22];

endmodule



module compressBy4_inWidth27
(
  in,
  out
);

  input [26:0] in;
  output [6:0] out;
  wire [6:0] out;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;
  assign out[0] = N1 | in[0];
  assign N1 = N0 | in[1];
  assign N0 = in[3] | in[2];
  assign out[1] = N3 | in[4];
  assign N3 = N2 | in[5];
  assign N2 = in[7] | in[6];
  assign out[2] = N5 | in[8];
  assign N5 = N4 | in[9];
  assign N4 = in[11] | in[10];
  assign out[3] = N7 | in[12];
  assign N7 = N6 | in[13];
  assign N6 = in[15] | in[14];
  assign out[4] = N9 | in[16];
  assign N9 = N8 | in[17];
  assign N8 = in[19] | in[18];
  assign out[5] = N11 | in[20];
  assign N11 = N10 | in[21];
  assign N10 = in[23] | in[22];
  assign out[6] = N12 | in[24];
  assign N12 = in[26] | in[25];

endmodule



module reverse_width6
(
  in,
  out
);

  input [5:0] in;
  output [5:0] out;
  wire [5:0] out;
  assign out[5] = in[0];
  assign out[4] = in[1];
  assign out[3] = in[2];
  assign out[2] = in[3];
  assign out[1] = in[4];
  assign out[0] = in[5];

endmodule



module lowMaskHiLo_inWidth5_topBound18_bottomBound12
(
  in,
  out
);

  input [4:0] in;
  output [5:0] out;
  wire [5:0] out,reverseOut;
  wire sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13;

  reverse_width6
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> in;

endmodule



module mulAddRecFNToRaw_preMul_8_24_1
(
  control,
  op,
  a,
  b,
  c,
  roundingMode,
  mulAddA,
  mulAddB,
  mulAddC,
  intermed_compactState,
  intermed_sExp,
  intermed_CDom_CAlignDist,
  intermed_highAlignedSigC
);

  input [0:0] control;
  input [2:0] op;
  input [32:0] a;
  input [32:0] b;
  input [32:0] c;
  input [2:0] roundingMode;
  output [23:0] mulAddA;
  output [23:0] mulAddB;
  output [47:0] mulAddC;
  output [5:0] intermed_compactState;
  output [9:0] intermed_sExp;
  output [4:0] intermed_CDom_CAlignDist;
  output [25:0] intermed_highAlignedSigC;
  wire [23:0] mulAddA,mulAddB;
  wire [47:0] mulAddC;
  wire [5:0] intermed_compactState,CExtraMask;
  wire [9:0] intermed_sExp,sExpA,sExpB,sExpC;
  wire [4:0] intermed_CDom_CAlignDist;
  wire [25:0] intermed_highAlignedSigC;
  wire N0,N1,N2,N3,N4,N5,isNaNA,isInfA,isZeroA,signA,isSigNaNA,isNaNB,isInfB,isZeroB,
  signB,isSigNaNB,isNaNC,isInfC,isZeroC,signC,isSigNaNC,signProd,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,opSignC,N17,isMinCAlign,N18,CIsDominant,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  reduced4CExtra,N61,N62,isNaNAOrB,isNaNAny,isInfAOrB,invalidProd,notSigNaN_invalidExc,
  invalidExc,notNaN_addZeros,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,sv2v_dc_1;
  wire [24:0] sigA,sigB,sigC;
  wire [10:0] sExpAlignedProd,sNatCAlignDist;
  wire [6:5] CAlignDist;
  wire [77:52] extComplSigC;
  wire [50:0] mainAlignedSigC;
  wire [6:0] reduced4SigC;
  wire [0:0] alignedSigC;
  wire [7:0] \fi1.aux_part ;

  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN_a
  (
    .in(a),
    .isNaN(isNaNA),
    .isInf(isInfA),
    .isZero(isZeroA),
    .sign(signA),
    .sExp(sExpA),
    .sig(sigA)
  );


  isSigNaNRecFN_expWidth8_sigWidth24
  isSigNaN_a
  (
    .in(a),
    .isSigNaN(isSigNaNA)
  );


  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN_b
  (
    .in(b),
    .isNaN(isNaNB),
    .isInf(isInfB),
    .isZero(isZeroB),
    .sign(signB),
    .sExp(sExpB),
    .sig(sigB)
  );


  isSigNaNRecFN_expWidth8_sigWidth24
  isSigNaN_b
  (
    .in(b),
    .isSigNaN(isSigNaNB)
  );


  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN_c
  (
    .in(c),
    .isNaN(isNaNC),
    .isInf(isInfC),
    .isZero(isZeroC),
    .sign(signC),
    .sExp(sExpC),
    .sig(sigC)
  );


  isSigNaNRecFN_expWidth8_sigWidth24
  isSigNaN_c
  (
    .in(c),
    .isSigNaN(isSigNaNC)
  );

  assign N17 = $signed(sNatCAlignDist) < $signed(1'b0);
  assign N18 = sNatCAlignDist[9:0] <= { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 };
  assign N30 = sNatCAlignDist[9:0] < { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 };
  assign { sv2v_dc_1, intermed_highAlignedSigC, mainAlignedSigC } = $signed({ extComplSigC, extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52], extComplSigC[52:52] }) >>> { CAlignDist, intermed_CDom_CAlignDist };

  compressBy4_inWidth27
  compressBy4_sigC
  (
    .in({ sigC, 1'b0, 1'b0 }),
    .out(reduced4SigC)
  );


  lowMaskHiLo_inWidth5_topBound18_bottomBound12
  lowMask_CExtraMask
  (
    .in({ CAlignDist, intermed_CDom_CAlignDist[4:2] }),
    .out(CExtraMask)
  );

  assign N80 = ~roundingMode[1];
  assign N81 = N80 | roundingMode[2];
  assign N82 = roundingMode[0] | N81;
  assign N83 = ~N82;
  assign { N71, N70, N69, N68, N67, N66, N65, N64 } = a[7:0] * b[31:24];
  assign { N79, N78, N77, N76, N75, N74, N73, N72 } = a[31:24] * b[7:0];
  assign { N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6 } = $signed(sExpA) + $signed(sExpB);
  assign \fi1.aux_part  = { N71, N70, N69, N68, N67, N66, N65, N64 } + { N79, N78, N77, N76, N75, N74, N73, N72 };
  assign sExpAlignedProd = $signed({ N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6 }) + $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 });
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(sExpC);
  assign { N29, N28, N27, N26, N25, N24, N23, N22, N21, N20 } = $signed(sExpAlignedProd[9:0]) - $signed({ 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 });
  assign intermed_sExp = (N0)? sExpC : 
                         (N1)? { N29, N28, N27, N26, N25, N24, N23, N22, N21, N20 } : 1'b0;
  assign N0 = CIsDominant;
  assign N1 = N19;
  assign { CAlignDist, intermed_CDom_CAlignDist } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                    (N34)? sNatCAlignDist[6:0] : 
                                                    (N32)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign N2 = isMinCAlign;
  assign extComplSigC[77:53] = (N3)? { N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60 } : 
                               (N4)? sigC : 1'b0;
  assign N3 = extComplSigC[52];
  assign N4 = N35;
  assign alignedSigC[0] = (N3)? N61 : 
                          (N4)? N62 : 1'b0;
  assign mulAddA = (N5)? a[23:0] : 
                   (N63)? sigA[23:0] : 1'b0;
  assign N5 = op[2];
  assign mulAddB = (N5)? b[23:0] : 
                   (N63)? sigB[23:0] : 1'b0;
  assign mulAddC = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \fi1.aux_part , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                   (N63)? mainAlignedSigC[50:3] : 1'b0;
  assign signProd = N84 ^ op[1];
  assign N84 = signA ^ signB;
  assign extComplSigC[52] = N85 ^ op[0];
  assign N85 = signProd ^ signC;
  assign opSignC = signProd ^ extComplSigC[52];
  assign isMinCAlign = N86 | N17;
  assign N86 = isZeroA | isZeroB;
  assign CIsDominant = N87 & N88;
  assign N87 = ~isZeroC;
  assign N88 = isMinCAlign | N18;
  assign N19 = ~CIsDominant;
  assign N31 = N30 | isMinCAlign;
  assign N32 = ~N31;
  assign N33 = ~isMinCAlign;
  assign N34 = N30 & N33;
  assign N35 = ~extComplSigC[52];
  assign N36 = ~sigC[24];
  assign N37 = ~sigC[23];
  assign N38 = ~sigC[22];
  assign N39 = ~sigC[21];
  assign N40 = ~sigC[20];
  assign N41 = ~sigC[19];
  assign N42 = ~sigC[18];
  assign N43 = ~sigC[17];
  assign N44 = ~sigC[16];
  assign N45 = ~sigC[15];
  assign N46 = ~sigC[14];
  assign N47 = ~sigC[13];
  assign N48 = ~sigC[12];
  assign N49 = ~sigC[11];
  assign N50 = ~sigC[10];
  assign N51 = ~sigC[9];
  assign N52 = ~sigC[8];
  assign N53 = ~sigC[7];
  assign N54 = ~sigC[6];
  assign N55 = ~sigC[5];
  assign N56 = ~sigC[4];
  assign N57 = ~sigC[3];
  assign N58 = ~sigC[2];
  assign N59 = ~sigC[1];
  assign N60 = ~sigC[0];
  assign reduced4CExtra = N97 | N98;
  assign N97 = N95 | N96;
  assign N95 = N93 | N94;
  assign N93 = N91 | N92;
  assign N91 = N89 | N90;
  assign N89 = reduced4SigC[5] & CExtraMask[5];
  assign N90 = reduced4SigC[4] & CExtraMask[4];
  assign N92 = reduced4SigC[3] & CExtraMask[3];
  assign N94 = reduced4SigC[2] & CExtraMask[2];
  assign N96 = reduced4SigC[1] & CExtraMask[1];
  assign N98 = reduced4SigC[0] & CExtraMask[0];
  assign N61 = N100 & N101;
  assign N100 = N99 & mainAlignedSigC[0];
  assign N99 = mainAlignedSigC[2] & mainAlignedSigC[1];
  assign N101 = ~reduced4CExtra;
  assign N62 = N103 | reduced4CExtra;
  assign N103 = N102 | mainAlignedSigC[0];
  assign N102 = mainAlignedSigC[2] | mainAlignedSigC[1];
  assign isNaNAOrB = isNaNA | isNaNB;
  assign isNaNAny = isNaNAOrB | isNaNC;
  assign isInfAOrB = isInfA | isInfB;
  assign invalidProd = N104 | N105;
  assign N104 = isInfA & isZeroB;
  assign N105 = isZeroA & isInfB;
  assign notSigNaN_invalidExc = invalidProd | N109;
  assign N109 = N108 & extComplSigC[52];
  assign N108 = N107 & isInfC;
  assign N107 = N106 & isInfAOrB;
  assign N106 = ~isNaNAOrB;
  assign invalidExc = N111 | notSigNaN_invalidExc;
  assign N111 = N110 | isSigNaNC;
  assign N110 = isSigNaNA | isSigNaNB;
  assign notNaN_addZeros = N112 & isZeroC;
  assign N112 = isZeroA | isZeroB;
  assign intermed_compactState[5] = N114 | notNaN_addZeros;
  assign N114 = N113 | isInfC;
  assign N113 = isNaNAny | isInfAOrB;
  assign intermed_compactState[0] = N121 | N124;
  assign N121 = N117 | N120;
  assign N117 = N115 | N116;
  assign N115 = isInfAOrB & signProd;
  assign N116 = isInfC & opSignC;
  assign N120 = N119 & opSignC;
  assign N119 = N118 & signProd;
  assign N118 = notNaN_addZeros & N82;
  assign N124 = N122 & N123;
  assign N122 = notNaN_addZeros & N83;
  assign N123 = signProd | opSignC;
  assign N63 = ~op[2];
  assign intermed_compactState[4] = invalidExc | N126;
  assign N126 = N125 & signProd;
  assign N125 = ~intermed_compactState[5];
  assign intermed_compactState[3] = isNaNAny | N127;
  assign N127 = N125 & extComplSigC[52];
  assign intermed_compactState[2] = N128 | N129;
  assign N128 = isInfAOrB | isInfC;
  assign N129 = N125 & CIsDominant;
  assign intermed_compactState[1] = notNaN_addZeros | N130;
  assign N130 = N125 & alignedSigC[0];

endmodule



module lowMaskLoHi_inWidth3_topBound0_bottomBound6
(
  in,
  out
);

  input [2:0] in;
  output [5:0] out;
  wire [5:0] out,reverseOut;
  wire N0,N1,N2,sv2v_dc_1,sv2v_dc_2;

  reverse_width6
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { N0, N1, N2 };
  assign N0 = ~in[2];
  assign N1 = ~in[1];
  assign N2 = ~in[0];

endmodule



module compressBy2_inWidth51
(
  in,
  out
);

  input [50:0] in;
  output [25:0] out;
  wire [25:0] out;
  wire out_25_;
  assign out_25_ = in[50];
  assign out[25] = out_25_;
  assign out[0] = in[1] | in[0];
  assign out[1] = in[3] | in[2];
  assign out[2] = in[5] | in[4];
  assign out[3] = in[7] | in[6];
  assign out[4] = in[9] | in[8];
  assign out[5] = in[11] | in[10];
  assign out[6] = in[13] | in[12];
  assign out[7] = in[15] | in[14];
  assign out[8] = in[17] | in[16];
  assign out[9] = in[19] | in[18];
  assign out[10] = in[21] | in[20];
  assign out[11] = in[23] | in[22];
  assign out[12] = in[25] | in[24];
  assign out[13] = in[27] | in[26];
  assign out[14] = in[29] | in[28];
  assign out[15] = in[31] | in[30];
  assign out[16] = in[33] | in[32];
  assign out[17] = in[35] | in[34];
  assign out[18] = in[37] | in[36];
  assign out[19] = in[39] | in[38];
  assign out[20] = in[41] | in[40];
  assign out[21] = in[43] | in[42];
  assign out[22] = in[45] | in[44];
  assign out[23] = in[47] | in[46];
  assign out[24] = in[49] | in[48];

endmodule



module reverse_width26
(
  in,
  out
);

  input [25:0] in;
  output [25:0] out;
  wire [25:0] out;
  assign out[25] = in[0];
  assign out[24] = in[1];
  assign out[23] = in[2];
  assign out[22] = in[3];
  assign out[21] = in[4];
  assign out[20] = in[5];
  assign out[19] = in[6];
  assign out[18] = in[7];
  assign out[17] = in[8];
  assign out[16] = in[9];
  assign out[15] = in[10];
  assign out[14] = in[11];
  assign out[13] = in[12];
  assign out[12] = in[13];
  assign out[11] = in[14];
  assign out[10] = in[15];
  assign out[9] = in[16];
  assign out[8] = in[17];
  assign out[7] = in[18];
  assign out[6] = in[19];
  assign out[5] = in[20];
  assign out[4] = in[21];
  assign out[3] = in[22];
  assign out[2] = in[23];
  assign out[1] = in[24];
  assign out[0] = in[25];

endmodule



module countLeadingZeros_inWidth26_countWidth5
(
  in,
  count
);

  input [25:0] in;
  output [4:0] count;
  wire [4:0] count;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,\Bit_5_.countSoFar_0 ,\Bit_9_.countSoFar_0 ,
  \Bit_10_.countSoFar_1 ,\Bit_11_.countSoFar_3 ,\Bit_13_.countSoFar_0 ,
  \Bit_17_.countSoFar_0 ,\Bit_18_.countSoFar_1 ,\Bit_19_.countSoFar_4 ,\Bit_20_.countSoFar_2 ,
  \Bit_21_.countSoFar_2 ,\Bit_21_.countSoFar_0 ,\Bit_22_.countSoFar_4 ,
  \Bit_23_.countSoFar_4 ,sv2v_dc_1;
  wire [25:0] reverseIn;
  wire [26:1] oneLeastReverseIn;
  wire [0:0] \Bit_1_.countSoFar ;
  wire [1:1] \Bit_2_.countSoFar ;
  wire [1:0] \Bit_3_.countSoFar ,\Bit_11_.countSoFar ,\Bit_19_.countSoFar ,
  \Bit_23_.countSoFar ;
  wire [2:2] \Bit_4_.countSoFar ,\Bit_5_.countSoFar ;
  wire [2:1] \Bit_6_.countSoFar ,\Bit_22_.countSoFar ;
  wire [2:0] \Bit_7_.countSoFar ;
  wire [3:3] \Bit_8_.countSoFar ,\Bit_9_.countSoFar ,\Bit_10_.countSoFar ;
  wire [3:2] \Bit_12_.countSoFar ,\Bit_13_.countSoFar ;
  wire [3:1] \Bit_14_.countSoFar ;
  wire [3:0] \Bit_15_.countSoFar ;
  wire [4:4] \Bit_16_.countSoFar ,\Bit_17_.countSoFar ,\Bit_18_.countSoFar ,
  \Bit_20_.countSoFar ,\Bit_21_.countSoFar ;
  wire [4:3] \Bit_24_.countSoFar ,\Bit_25_.countSoFar ;

  reverse_width26
  reverse_in
  (
    .in(in),
    .out(reverseIn)
  );

  assign { oneLeastReverseIn[26:26], N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, sv2v_dc_1 } = { N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25 } + 1'b1;
  assign N0 = ~reverseIn[25];
  assign N1 = ~reverseIn[24];
  assign N2 = ~reverseIn[23];
  assign N3 = ~reverseIn[22];
  assign N4 = ~reverseIn[21];
  assign N5 = ~reverseIn[20];
  assign N6 = ~reverseIn[19];
  assign N7 = ~reverseIn[18];
  assign N8 = ~reverseIn[17];
  assign N9 = ~reverseIn[16];
  assign N10 = ~reverseIn[15];
  assign N11 = ~reverseIn[14];
  assign N12 = ~reverseIn[13];
  assign N13 = ~reverseIn[12];
  assign N14 = ~reverseIn[11];
  assign N15 = ~reverseIn[10];
  assign N16 = ~reverseIn[9];
  assign N17 = ~reverseIn[8];
  assign N18 = ~reverseIn[7];
  assign N19 = ~reverseIn[6];
  assign N20 = ~reverseIn[5];
  assign N21 = ~reverseIn[4];
  assign N22 = ~reverseIn[3];
  assign N23 = ~reverseIn[2];
  assign N24 = ~reverseIn[1];
  assign N25 = ~reverseIn[0];
  assign oneLeastReverseIn[25] = reverseIn[25] & N50;
  assign oneLeastReverseIn[24] = reverseIn[24] & N49;
  assign oneLeastReverseIn[23] = reverseIn[23] & N48;
  assign oneLeastReverseIn[22] = reverseIn[22] & N47;
  assign oneLeastReverseIn[21] = reverseIn[21] & N46;
  assign oneLeastReverseIn[20] = reverseIn[20] & N45;
  assign oneLeastReverseIn[19] = reverseIn[19] & N44;
  assign oneLeastReverseIn[18] = reverseIn[18] & N43;
  assign oneLeastReverseIn[17] = reverseIn[17] & N42;
  assign oneLeastReverseIn[16] = reverseIn[16] & N41;
  assign oneLeastReverseIn[15] = reverseIn[15] & N40;
  assign oneLeastReverseIn[14] = reverseIn[14] & N39;
  assign oneLeastReverseIn[13] = reverseIn[13] & N38;
  assign oneLeastReverseIn[12] = reverseIn[12] & N37;
  assign oneLeastReverseIn[11] = reverseIn[11] & N36;
  assign oneLeastReverseIn[10] = reverseIn[10] & N35;
  assign oneLeastReverseIn[9] = reverseIn[9] & N34;
  assign oneLeastReverseIn[8] = reverseIn[8] & N33;
  assign oneLeastReverseIn[7] = reverseIn[7] & N32;
  assign oneLeastReverseIn[6] = reverseIn[6] & N31;
  assign oneLeastReverseIn[5] = reverseIn[5] & N30;
  assign oneLeastReverseIn[4] = reverseIn[4] & N29;
  assign oneLeastReverseIn[3] = reverseIn[3] & N28;
  assign oneLeastReverseIn[2] = reverseIn[2] & N27;
  assign oneLeastReverseIn[1] = reverseIn[1] & N26;
  assign \Bit_1_.countSoFar [0] = 1'b0 | oneLeastReverseIn[1];
  assign \Bit_2_.countSoFar [1] = 1'b0 | oneLeastReverseIn[2];
  assign \Bit_3_.countSoFar [1] = \Bit_2_.countSoFar [1] | oneLeastReverseIn[3];
  assign \Bit_3_.countSoFar [0] = \Bit_1_.countSoFar [0] | oneLeastReverseIn[3];
  assign \Bit_4_.countSoFar [2] = 1'b0 | oneLeastReverseIn[4];
  assign \Bit_5_.countSoFar [2] = \Bit_4_.countSoFar [2] | oneLeastReverseIn[5];
  assign \Bit_5_.countSoFar_0  = \Bit_3_.countSoFar [0] | oneLeastReverseIn[5];
  assign \Bit_6_.countSoFar [2] = \Bit_5_.countSoFar [2] | oneLeastReverseIn[6];
  assign \Bit_6_.countSoFar [1] = \Bit_3_.countSoFar [1] | oneLeastReverseIn[6];
  assign \Bit_7_.countSoFar [2] = \Bit_6_.countSoFar [2] | oneLeastReverseIn[7];
  assign \Bit_7_.countSoFar [1] = \Bit_6_.countSoFar [1] | oneLeastReverseIn[7];
  assign \Bit_7_.countSoFar [0] = \Bit_5_.countSoFar_0  | oneLeastReverseIn[7];
  assign \Bit_8_.countSoFar [3] = 1'b0 | oneLeastReverseIn[8];
  assign \Bit_9_.countSoFar [3] = \Bit_8_.countSoFar [3] | oneLeastReverseIn[9];
  assign \Bit_9_.countSoFar_0  = \Bit_7_.countSoFar [0] | oneLeastReverseIn[9];
  assign \Bit_10_.countSoFar [3] = \Bit_9_.countSoFar [3] | oneLeastReverseIn[10];
  assign \Bit_10_.countSoFar_1  = \Bit_7_.countSoFar [1] | oneLeastReverseIn[10];
  assign \Bit_11_.countSoFar_3  = \Bit_10_.countSoFar [3] | oneLeastReverseIn[11];
  assign \Bit_11_.countSoFar [1] = \Bit_10_.countSoFar_1  | oneLeastReverseIn[11];
  assign \Bit_11_.countSoFar [0] = \Bit_9_.countSoFar_0  | oneLeastReverseIn[11];
  assign \Bit_12_.countSoFar [3] = \Bit_11_.countSoFar_3  | oneLeastReverseIn[12];
  assign \Bit_12_.countSoFar [2] = \Bit_7_.countSoFar [2] | oneLeastReverseIn[12];
  assign \Bit_13_.countSoFar [3] = \Bit_12_.countSoFar [3] | oneLeastReverseIn[13];
  assign \Bit_13_.countSoFar [2] = \Bit_12_.countSoFar [2] | oneLeastReverseIn[13];
  assign \Bit_13_.countSoFar_0  = \Bit_11_.countSoFar [0] | oneLeastReverseIn[13];
  assign \Bit_14_.countSoFar [3] = \Bit_13_.countSoFar [3] | oneLeastReverseIn[14];
  assign \Bit_14_.countSoFar [2] = \Bit_13_.countSoFar [2] | oneLeastReverseIn[14];
  assign \Bit_14_.countSoFar [1] = \Bit_11_.countSoFar [1] | oneLeastReverseIn[14];
  assign \Bit_15_.countSoFar [3] = \Bit_14_.countSoFar [3] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [2] = \Bit_14_.countSoFar [2] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [1] = \Bit_14_.countSoFar [1] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [0] = \Bit_13_.countSoFar_0  | oneLeastReverseIn[15];
  assign \Bit_16_.countSoFar [4] = 1'b0 | oneLeastReverseIn[16];
  assign \Bit_17_.countSoFar [4] = \Bit_16_.countSoFar [4] | oneLeastReverseIn[17];
  assign \Bit_17_.countSoFar_0  = \Bit_15_.countSoFar [0] | oneLeastReverseIn[17];
  assign \Bit_18_.countSoFar [4] = \Bit_17_.countSoFar [4] | oneLeastReverseIn[18];
  assign \Bit_18_.countSoFar_1  = \Bit_15_.countSoFar [1] | oneLeastReverseIn[18];
  assign \Bit_19_.countSoFar_4  = \Bit_18_.countSoFar [4] | oneLeastReverseIn[19];
  assign \Bit_19_.countSoFar [1] = \Bit_18_.countSoFar_1  | oneLeastReverseIn[19];
  assign \Bit_19_.countSoFar [0] = \Bit_17_.countSoFar_0  | oneLeastReverseIn[19];
  assign \Bit_20_.countSoFar [4] = \Bit_19_.countSoFar_4  | oneLeastReverseIn[20];
  assign \Bit_20_.countSoFar_2  = \Bit_15_.countSoFar [2] | oneLeastReverseIn[20];
  assign \Bit_21_.countSoFar [4] = \Bit_20_.countSoFar [4] | oneLeastReverseIn[21];
  assign \Bit_21_.countSoFar_2  = \Bit_20_.countSoFar_2  | oneLeastReverseIn[21];
  assign \Bit_21_.countSoFar_0  = \Bit_19_.countSoFar [0] | oneLeastReverseIn[21];
  assign \Bit_22_.countSoFar_4  = \Bit_21_.countSoFar [4] | oneLeastReverseIn[22];
  assign \Bit_22_.countSoFar [2] = \Bit_21_.countSoFar_2  | oneLeastReverseIn[22];
  assign \Bit_22_.countSoFar [1] = \Bit_19_.countSoFar [1] | oneLeastReverseIn[22];
  assign \Bit_23_.countSoFar_4  = \Bit_22_.countSoFar_4  | oneLeastReverseIn[23];
  assign count[2] = \Bit_22_.countSoFar [2] | oneLeastReverseIn[23];
  assign \Bit_23_.countSoFar [1] = \Bit_22_.countSoFar [1] | oneLeastReverseIn[23];
  assign \Bit_23_.countSoFar [0] = \Bit_21_.countSoFar_0  | oneLeastReverseIn[23];
  assign \Bit_24_.countSoFar [4] = \Bit_23_.countSoFar_4  | oneLeastReverseIn[24];
  assign \Bit_24_.countSoFar [3] = \Bit_15_.countSoFar [3] | oneLeastReverseIn[24];
  assign \Bit_25_.countSoFar [4] = \Bit_24_.countSoFar [4] | oneLeastReverseIn[25];
  assign \Bit_25_.countSoFar [3] = \Bit_24_.countSoFar [3] | oneLeastReverseIn[25];
  assign count[0] = \Bit_23_.countSoFar [0] | oneLeastReverseIn[25];
  assign count[4] = \Bit_25_.countSoFar [4] | oneLeastReverseIn[26];
  assign count[3] = \Bit_25_.countSoFar [3] | oneLeastReverseIn[26];
  assign count[1] = \Bit_23_.countSoFar [1] | oneLeastReverseIn[26];

endmodule



module compressBy2_inWidth13
(
  in,
  out
);

  input [12:0] in;
  output [6:0] out;
  wire [6:0] out;
  wire out_6_;
  assign out_6_ = in[12];
  assign out[6] = out_6_;
  assign out[0] = in[1] | in[0];
  assign out[1] = in[3] | in[2];
  assign out[2] = in[5] | in[4];
  assign out[3] = in[7] | in[6];
  assign out[4] = in[9] | in[8];
  assign out[5] = in[11] | in[10];

endmodule



module lowMaskLoHi_inWidth4_topBound0_bottomBound6
(
  in,
  out
);

  input [3:0] in;
  output [5:0] out;
  wire [5:0] out,reverseOut;
  wire N0,N1,N2,N3,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,
  sv2v_dc_7,sv2v_dc_8,sv2v_dc_9,sv2v_dc_10;

  reverse_width6
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { N0, N1, N2, N3 };
  assign N0 = ~in[3];
  assign N1 = ~in[2];
  assign N2 = ~in[1];
  assign N3 = ~in[0];

endmodule



module mulAddRecFNToRaw_postMul_expWidth8_sigWidth24
(
  intermed_compactState,
  intermed_sExp,
  intermed_CDom_CAlignDist,
  intermed_highAlignedSigC,
  mulAddResult,
  roundingMode,
  invalidExc,
  out_isNaN,
  out_isInf,
  out_isZero,
  out_sign,
  out_sExp,
  out_sig
);

  input [5:0] intermed_compactState;
  input [9:0] intermed_sExp;
  input [4:0] intermed_CDom_CAlignDist;
  input [25:0] intermed_highAlignedSigC;
  input [48:0] mulAddResult;
  input [2:0] roundingMode;
  output [9:0] out_sExp;
  output [26:0] out_sig;
  output invalidExc;
  output out_isNaN;
  output out_isInf;
  output out_isZero;
  output out_sign;
  wire [9:0] out_sExp,CDom_sExp,notCDom_sExp;
  wire [26:0] out_sig;
  wire invalidExc,out_isNaN,out_isInf,out_isZero,out_sign,N0,N1,N2,N3,N4,N5,N6,N7,N8,
  notNaN_addZeros,opSignC,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  CDom_absSigSumExtra,N62,CDom_reduced4SigExtra,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  notCDom_reduced4SigExtra,notCDom_completeCancellation,N139,notCDom_sign,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,
  sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,sv2v_dc_28,sv2v_dc_29,sv2v_dc_30,
  sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,
  sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,sv2v_dc_43,sv2v_dc_44;
  wire [25:0] incHighAlignedSigC,notCDom_reduced2AbsSigSum;
  wire [74:49] sigSum;
  wire [49:0] CDom_absSigSum;
  wire [28:0] CDom_mainSig,notCDom_mainSig;
  wire [6:0] CDom_reduced4LowSig,notCDom_reduced4AbsSigSum;
  wire [5:0] CDom_sigExtraMask,notCDom_sigExtraMask;
  wire [0:0] CDom_sig,notCDom_sig;
  wire [50:0] notCDom_absSigSum;
  wire [4:0] notCDom_normDistReduced2;
  assign { CDom_mainSig, sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21 } = CDom_absSigSum << intermed_CDom_CAlignDist;

  compressBy4_inWidth27
  compressBy4_CDom_absSigSum
  (
    .in({ CDom_absSigSum[23:0], 1'b0, 1'b0, 1'b0 }),
    .out(CDom_reduced4LowSig)
  );


  lowMaskLoHi_inWidth3_topBound0_bottomBound6
  lowMask_CDom_sigExtraMask
  (
    .in(intermed_CDom_CAlignDist[4:2]),
    .out(CDom_sigExtraMask)
  );


  compressBy2_inWidth51
  compressBy2_notCDom_absSigSum
  (
    .in(notCDom_absSigSum),
    .out(notCDom_reduced2AbsSigSum)
  );


  countLeadingZeros_inWidth26_countWidth5
  countLeadingZeros_notCDom
  (
    .in(notCDom_reduced2AbsSigSum),
    .count(notCDom_normDistReduced2)
  );

  assign { notCDom_mainSig, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44 } = { 1'b0, notCDom_absSigSum } << { notCDom_normDistReduced2, 1'b0 };

  compressBy2_inWidth13
  compressBy2_notCDom_reduced2AbsSigSum
  (
    .in(notCDom_reduced2AbsSigSum[12:0]),
    .out(notCDom_reduced4AbsSigSum)
  );


  lowMaskLoHi_inWidth4_topBound0_bottomBound6
  lowMask_notCDom_sigExtraMask
  (
    .in(notCDom_normDistReduced2[4:1]),
    .out(notCDom_sigExtraMask)
  );

  assign notCDom_completeCancellation = notCDom_mainSig[28:27] == 1'b0;
  assign N141 = ~roundingMode[1];
  assign N142 = N141 | roundingMode[2];
  assign N143 = roundingMode[0] | N142;
  assign N144 = ~N143;
  assign CDom_sExp = intermed_sExp - intermed_compactState[3];
  assign notCDom_sExp = intermed_sExp - { notCDom_normDistReduced2, 1'b0 };
  assign incHighAlignedSigC = intermed_highAlignedSigC + 1'b1;
  assign { N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88 } = { sigSum[50:49], mulAddResult[47:0], intermed_compactState[1:1] } + intermed_compactState[3];
  assign sigSum = (N0)? incHighAlignedSigC : 
                  (N9)? intermed_highAlignedSigC : 1'b0;
  assign N0 = mulAddResult[48];
  assign CDom_absSigSum = (N1)? { N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59 } : 
                          (N2)? { 1'b0, intermed_highAlignedSigC[25:24], sigSum[72:49], mulAddResult[47:25] } : 1'b0;
  assign N1 = intermed_compactState[3];
  assign N2 = N60;
  assign CDom_absSigSumExtra = (N1)? N61 : 
                               (N2)? N62 : 1'b0;
  assign notCDom_absSigSum = (N3)? { N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87 } : 
                             (N4)? { N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88 } : 1'b0;
  assign N3 = sigSum[51];
  assign N4 = N33;
  assign notCDom_sign = (N5)? N144 : 
                        (N6)? N140 : 1'b0;
  assign N5 = notCDom_completeCancellation;
  assign N6 = N139;
  assign out_sExp = (N7)? CDom_sExp : 
                    (N8)? notCDom_sExp : 1'b0;
  assign N7 = intermed_compactState[2];
  assign N8 = N216;
  assign out_sig = (N7)? { CDom_mainSig[28:3], CDom_sig[0:0] } : 
                   (N8)? { notCDom_mainSig[28:3], notCDom_sig[0:0] } : 1'b0;
  assign invalidExc = intermed_compactState[5] & intermed_compactState[4];
  assign out_isNaN = intermed_compactState[5] & intermed_compactState[3];
  assign out_isInf = intermed_compactState[5] & intermed_compactState[2];
  assign notNaN_addZeros = intermed_compactState[5] & intermed_compactState[1];
  assign opSignC = intermed_compactState[4] ^ intermed_compactState[3];
  assign N9 = ~mulAddResult[48];
  assign N10 = ~sigSum[74];
  assign N11 = ~sigSum[73];
  assign N12 = ~sigSum[72];
  assign N13 = ~sigSum[71];
  assign N14 = ~sigSum[70];
  assign N15 = ~sigSum[69];
  assign N16 = ~sigSum[68];
  assign N17 = ~sigSum[67];
  assign N18 = ~sigSum[66];
  assign N19 = ~sigSum[65];
  assign N20 = ~sigSum[64];
  assign N21 = ~sigSum[63];
  assign N22 = ~sigSum[62];
  assign N23 = ~sigSum[61];
  assign N24 = ~sigSum[60];
  assign N25 = ~sigSum[59];
  assign N26 = ~sigSum[58];
  assign N27 = ~sigSum[57];
  assign N28 = ~sigSum[56];
  assign N29 = ~sigSum[55];
  assign N30 = ~sigSum[54];
  assign N31 = ~sigSum[53];
  assign N32 = ~sigSum[52];
  assign N33 = ~sigSum[51];
  assign N34 = ~sigSum[50];
  assign N35 = ~sigSum[49];
  assign N36 = ~mulAddResult[47];
  assign N37 = ~mulAddResult[46];
  assign N38 = ~mulAddResult[45];
  assign N39 = ~mulAddResult[44];
  assign N40 = ~mulAddResult[43];
  assign N41 = ~mulAddResult[42];
  assign N42 = ~mulAddResult[41];
  assign N43 = ~mulAddResult[40];
  assign N44 = ~mulAddResult[39];
  assign N45 = ~mulAddResult[38];
  assign N46 = ~mulAddResult[37];
  assign N47 = ~mulAddResult[36];
  assign N48 = ~mulAddResult[35];
  assign N49 = ~mulAddResult[34];
  assign N50 = ~mulAddResult[33];
  assign N51 = ~mulAddResult[32];
  assign N52 = ~mulAddResult[31];
  assign N53 = ~mulAddResult[30];
  assign N54 = ~mulAddResult[29];
  assign N55 = ~mulAddResult[28];
  assign N56 = ~mulAddResult[27];
  assign N57 = ~mulAddResult[26];
  assign N58 = ~mulAddResult[25];
  assign N59 = ~mulAddResult[24];
  assign N60 = ~intermed_compactState[3];
  assign N61 = ~N167;
  assign N167 = N166 & mulAddResult[0];
  assign N166 = N165 & mulAddResult[1];
  assign N165 = N164 & mulAddResult[2];
  assign N164 = N163 & mulAddResult[3];
  assign N163 = N162 & mulAddResult[4];
  assign N162 = N161 & mulAddResult[5];
  assign N161 = N160 & mulAddResult[6];
  assign N160 = N159 & mulAddResult[7];
  assign N159 = N158 & mulAddResult[8];
  assign N158 = N157 & mulAddResult[9];
  assign N157 = N156 & mulAddResult[10];
  assign N156 = N155 & mulAddResult[11];
  assign N155 = N154 & mulAddResult[12];
  assign N154 = N153 & mulAddResult[13];
  assign N153 = N152 & mulAddResult[14];
  assign N152 = N151 & mulAddResult[15];
  assign N151 = N150 & mulAddResult[16];
  assign N150 = N149 & mulAddResult[17];
  assign N149 = N148 & mulAddResult[18];
  assign N148 = N147 & mulAddResult[19];
  assign N147 = N146 & mulAddResult[20];
  assign N146 = N145 & mulAddResult[21];
  assign N145 = mulAddResult[23] & mulAddResult[22];
  assign N62 = N190 | mulAddResult[0];
  assign N190 = N189 | mulAddResult[1];
  assign N189 = N188 | mulAddResult[2];
  assign N188 = N187 | mulAddResult[3];
  assign N187 = N186 | mulAddResult[4];
  assign N186 = N185 | mulAddResult[5];
  assign N185 = N184 | mulAddResult[6];
  assign N184 = N183 | mulAddResult[7];
  assign N183 = N182 | mulAddResult[8];
  assign N182 = N181 | mulAddResult[9];
  assign N181 = N180 | mulAddResult[10];
  assign N180 = N179 | mulAddResult[11];
  assign N179 = N178 | mulAddResult[12];
  assign N178 = N177 | mulAddResult[13];
  assign N177 = N176 | mulAddResult[14];
  assign N176 = N175 | mulAddResult[15];
  assign N175 = N174 | mulAddResult[16];
  assign N174 = N173 | mulAddResult[17];
  assign N173 = N172 | mulAddResult[18];
  assign N172 = N171 | mulAddResult[19];
  assign N171 = N170 | mulAddResult[20];
  assign N170 = N169 | mulAddResult[21];
  assign N169 = N168 | mulAddResult[22];
  assign N168 = mulAddResult[24] | mulAddResult[23];
  assign CDom_reduced4SigExtra = N199 | N200;
  assign N199 = N197 | N198;
  assign N197 = N195 | N196;
  assign N195 = N193 | N194;
  assign N193 = N191 | N192;
  assign N191 = CDom_reduced4LowSig[5] & CDom_sigExtraMask[5];
  assign N192 = CDom_reduced4LowSig[4] & CDom_sigExtraMask[4];
  assign N194 = CDom_reduced4LowSig[3] & CDom_sigExtraMask[3];
  assign N196 = CDom_reduced4LowSig[2] & CDom_sigExtraMask[2];
  assign N198 = CDom_reduced4LowSig[1] & CDom_sigExtraMask[1];
  assign N200 = CDom_reduced4LowSig[0] & CDom_sigExtraMask[0];
  assign CDom_sig[0] = N203 | CDom_absSigSumExtra;
  assign N203 = N202 | CDom_reduced4SigExtra;
  assign N202 = N201 | CDom_mainSig[0];
  assign N201 = CDom_mainSig[2] | CDom_mainSig[1];
  assign N63 = ~mulAddResult[23];
  assign N64 = ~mulAddResult[22];
  assign N65 = ~mulAddResult[21];
  assign N66 = ~mulAddResult[20];
  assign N67 = ~mulAddResult[19];
  assign N68 = ~mulAddResult[18];
  assign N69 = ~mulAddResult[17];
  assign N70 = ~mulAddResult[16];
  assign N71 = ~mulAddResult[15];
  assign N72 = ~mulAddResult[14];
  assign N73 = ~mulAddResult[13];
  assign N74 = ~mulAddResult[12];
  assign N75 = ~mulAddResult[11];
  assign N76 = ~mulAddResult[10];
  assign N77 = ~mulAddResult[9];
  assign N78 = ~mulAddResult[8];
  assign N79 = ~mulAddResult[7];
  assign N80 = ~mulAddResult[6];
  assign N81 = ~mulAddResult[5];
  assign N82 = ~mulAddResult[4];
  assign N83 = ~mulAddResult[3];
  assign N84 = ~mulAddResult[2];
  assign N85 = ~mulAddResult[1];
  assign N86 = ~mulAddResult[0];
  assign N87 = ~intermed_compactState[1];
  assign notCDom_reduced4SigExtra = N212 | N213;
  assign N212 = N210 | N211;
  assign N210 = N208 | N209;
  assign N208 = N206 | N207;
  assign N206 = N204 | N205;
  assign N204 = notCDom_reduced4AbsSigSum[5] & notCDom_sigExtraMask[5];
  assign N205 = notCDom_reduced4AbsSigSum[4] & notCDom_sigExtraMask[4];
  assign N207 = notCDom_reduced4AbsSigSum[3] & notCDom_sigExtraMask[3];
  assign N209 = notCDom_reduced4AbsSigSum[2] & notCDom_sigExtraMask[2];
  assign N211 = notCDom_reduced4AbsSigSum[1] & notCDom_sigExtraMask[1];
  assign N213 = notCDom_reduced4AbsSigSum[0] & notCDom_sigExtraMask[0];
  assign notCDom_sig[0] = N215 | notCDom_reduced4SigExtra;
  assign N215 = N214 | notCDom_mainSig[0];
  assign N214 = notCDom_mainSig[2] | notCDom_mainSig[1];
  assign N139 = ~notCDom_completeCancellation;
  assign N140 = intermed_compactState[4] ^ sigSum[51];
  assign out_isZero = notNaN_addZeros | N217;
  assign N217 = N216 & notCDom_completeCancellation;
  assign N216 = ~intermed_compactState[2];
  assign out_sign = N222 | N224;
  assign N222 = N218 | N221;
  assign N218 = intermed_compactState[5] & intermed_compactState[0];
  assign N221 = N220 & opSignC;
  assign N220 = N219 & intermed_compactState[2];
  assign N219 = ~intermed_compactState[5];
  assign N224 = N223 & notCDom_sign;
  assign N223 = N219 & N216;

endmodule



module mulAddRecFNToRaw_expWidth8_sigWidth24
(
  control,
  op,
  a,
  b,
  c,
  roundingMode,
  invalidExc,
  out_isNaN,
  out_isInf,
  out_isZero,
  out_sign,
  out_sExp,
  out_sig,
  out_imul
);

  input [0:0] control;
  input [2:0] op;
  input [32:0] a;
  input [32:0] b;
  input [32:0] c;
  input [2:0] roundingMode;
  output [9:0] out_sExp;
  output [26:0] out_sig;
  output [31:0] out_imul;
  output invalidExc;
  output out_isNaN;
  output out_isInf;
  output out_isZero;
  output out_sign;
  wire [9:0] out_sExp,intermed_sExp;
  wire [26:0] out_sig;
  wire [31:0] out_imul;
  wire invalidExc,out_isNaN,out_isInf,out_isZero,out_sign,N0,N1,N2,N3,N4,N5,N6,N7,N8,
  N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,
  N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47;
  wire [23:0] mulAddA,mulAddB;
  wire [47:0] mulAddC;
  wire [5:0] intermed_compactState;
  wire [4:0] intermed_CDom_CAlignDist;
  wire [25:0] intermed_highAlignedSigC;
  wire [48:32] mulAddResult;

  mulAddRecFNToRaw_preMul_8_24_1
  mulAddToRaw_preMul
  (
    .control(control[0]),
    .op(op),
    .a(a),
    .b(b),
    .c(c),
    .roundingMode(roundingMode),
    .mulAddA(mulAddA),
    .mulAddB(mulAddB),
    .mulAddC(mulAddC),
    .intermed_compactState(intermed_compactState),
    .intermed_sExp(intermed_sExp),
    .intermed_CDom_CAlignDist(intermed_CDom_CAlignDist),
    .intermed_highAlignedSigC(intermed_highAlignedSigC)
  );


  mulAddRecFNToRaw_postMul_expWidth8_sigWidth24
  mulAddToRaw_postMul
  (
    .intermed_compactState(intermed_compactState),
    .intermed_sExp(intermed_sExp),
    .intermed_CDom_CAlignDist(intermed_CDom_CAlignDist),
    .intermed_highAlignedSigC(intermed_highAlignedSigC),
    .mulAddResult({ mulAddResult, out_imul }),
    .roundingMode(roundingMode),
    .invalidExc(invalidExc),
    .out_isNaN(out_isNaN),
    .out_isInf(out_isInf),
    .out_isZero(out_isZero),
    .out_sign(out_sign),
    .out_sExp(out_sExp),
    .out_sig(out_sig)
  );

  assign { N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } = mulAddA * mulAddB;
  assign { mulAddResult, out_imul } = { N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0 } + mulAddC;

endmodule



module fpu_float_fma
(
  clk_i,
  reset_i,
  stall_fpu1_i,
  imul_v_i,
  imul_rs1_i,
  imul_rs2_i,
  fp_v_i,
  fpu_float_op_i,
  fp_rs1_i,
  fp_rs2_i,
  fp_rs3_i,
  fp_rm_i,
  imul_v_o,
  imul_result_o,
  fma1_v_o,
  fma1_rm_o,
  invalidExc_o,
  out_isNaN_o,
  out_isInf_o,
  out_isZero_o,
  out_sign_o,
  out_sExp_o,
  out_sig_o
);

  input [31:0] imul_rs1_i;
  input [31:0] imul_rs2_i;
  input [3:0] fpu_float_op_i;
  input [32:0] fp_rs1_i;
  input [32:0] fp_rs2_i;
  input [32:0] fp_rs3_i;
  input [2:0] fp_rm_i;
  output [31:0] imul_result_o;
  output [2:0] fma1_rm_o;
  output [9:0] out_sExp_o;
  output [26:0] out_sig_o;
  input clk_i;
  input reset_i;
  input stall_fpu1_i;
  input imul_v_i;
  input fp_v_i;
  output imul_v_o;
  output fma1_v_o;
  output invalidExc_o;
  output out_isNaN_o;
  output out_isInf_o;
  output out_isZero_o;
  output out_sign_o;
  wire [31:0] imul_result_o,out_imul;
  wire [2:0] fma1_rm_o,fma_op_li;
  wire [9:0] out_sExp_o,out_sExp;
  wire [26:0] out_sig_o,out_sig;
  wire imul_v_o,fma1_v_o,invalidExc_o,out_isNaN_o,out_isInf_o,out_isZero_o,out_sign_o,
  N0,N1,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,is_fma_op,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,invalidExc,out_isNaN,out_isInf,out_isZero,out_sign,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132;
  wire [32:0] fma_a_li,fma_b_li,fma_c_li;
  reg imul_result_o_31_sv2v_reg,imul_result_o_30_sv2v_reg,imul_result_o_29_sv2v_reg,
  imul_result_o_28_sv2v_reg,imul_result_o_27_sv2v_reg,imul_result_o_26_sv2v_reg,
  imul_result_o_25_sv2v_reg,imul_result_o_24_sv2v_reg,imul_result_o_23_sv2v_reg,
  imul_result_o_22_sv2v_reg,imul_result_o_21_sv2v_reg,imul_result_o_20_sv2v_reg,
  imul_result_o_19_sv2v_reg,imul_result_o_18_sv2v_reg,imul_result_o_17_sv2v_reg,
  imul_result_o_16_sv2v_reg,imul_result_o_15_sv2v_reg,imul_result_o_14_sv2v_reg,
  imul_result_o_13_sv2v_reg,imul_result_o_12_sv2v_reg,imul_result_o_11_sv2v_reg,
  imul_result_o_10_sv2v_reg,imul_result_o_9_sv2v_reg,imul_result_o_8_sv2v_reg,
  imul_result_o_7_sv2v_reg,imul_result_o_6_sv2v_reg,imul_result_o_5_sv2v_reg,
  imul_result_o_4_sv2v_reg,imul_result_o_3_sv2v_reg,imul_result_o_2_sv2v_reg,imul_result_o_1_sv2v_reg,
  imul_result_o_0_sv2v_reg,fma1_v_o_sv2v_reg,fma1_rm_o_2_sv2v_reg,
  fma1_rm_o_1_sv2v_reg,fma1_rm_o_0_sv2v_reg,imul_v_o_sv2v_reg,out_sig_o_26_sv2v_reg,
  out_sig_o_25_sv2v_reg,out_sig_o_24_sv2v_reg,out_sig_o_23_sv2v_reg,out_sig_o_22_sv2v_reg,
  out_sig_o_21_sv2v_reg,out_sig_o_20_sv2v_reg,out_sig_o_19_sv2v_reg,out_sig_o_18_sv2v_reg,
  out_sig_o_17_sv2v_reg,out_sig_o_16_sv2v_reg,out_sig_o_15_sv2v_reg,
  out_sig_o_14_sv2v_reg,out_sig_o_13_sv2v_reg,out_sig_o_12_sv2v_reg,out_sig_o_11_sv2v_reg,
  out_sig_o_10_sv2v_reg,out_sig_o_9_sv2v_reg,out_sig_o_8_sv2v_reg,out_sig_o_7_sv2v_reg,
  out_sig_o_6_sv2v_reg,out_sig_o_5_sv2v_reg,out_sig_o_4_sv2v_reg,
  out_sig_o_3_sv2v_reg,out_sig_o_2_sv2v_reg,out_sig_o_1_sv2v_reg,out_sig_o_0_sv2v_reg,
  invalidExc_o_sv2v_reg,out_isNaN_o_sv2v_reg,out_isInf_o_sv2v_reg,out_isZero_o_sv2v_reg,
  out_sign_o_sv2v_reg,out_sExp_o_9_sv2v_reg,out_sExp_o_8_sv2v_reg,out_sExp_o_7_sv2v_reg,
  out_sExp_o_6_sv2v_reg,out_sExp_o_5_sv2v_reg,out_sExp_o_4_sv2v_reg,
  out_sExp_o_3_sv2v_reg,out_sExp_o_2_sv2v_reg,out_sExp_o_1_sv2v_reg,out_sExp_o_0_sv2v_reg;
  assign imul_result_o[31] = imul_result_o_31_sv2v_reg;
  assign imul_result_o[30] = imul_result_o_30_sv2v_reg;
  assign imul_result_o[29] = imul_result_o_29_sv2v_reg;
  assign imul_result_o[28] = imul_result_o_28_sv2v_reg;
  assign imul_result_o[27] = imul_result_o_27_sv2v_reg;
  assign imul_result_o[26] = imul_result_o_26_sv2v_reg;
  assign imul_result_o[25] = imul_result_o_25_sv2v_reg;
  assign imul_result_o[24] = imul_result_o_24_sv2v_reg;
  assign imul_result_o[23] = imul_result_o_23_sv2v_reg;
  assign imul_result_o[22] = imul_result_o_22_sv2v_reg;
  assign imul_result_o[21] = imul_result_o_21_sv2v_reg;
  assign imul_result_o[20] = imul_result_o_20_sv2v_reg;
  assign imul_result_o[19] = imul_result_o_19_sv2v_reg;
  assign imul_result_o[18] = imul_result_o_18_sv2v_reg;
  assign imul_result_o[17] = imul_result_o_17_sv2v_reg;
  assign imul_result_o[16] = imul_result_o_16_sv2v_reg;
  assign imul_result_o[15] = imul_result_o_15_sv2v_reg;
  assign imul_result_o[14] = imul_result_o_14_sv2v_reg;
  assign imul_result_o[13] = imul_result_o_13_sv2v_reg;
  assign imul_result_o[12] = imul_result_o_12_sv2v_reg;
  assign imul_result_o[11] = imul_result_o_11_sv2v_reg;
  assign imul_result_o[10] = imul_result_o_10_sv2v_reg;
  assign imul_result_o[9] = imul_result_o_9_sv2v_reg;
  assign imul_result_o[8] = imul_result_o_8_sv2v_reg;
  assign imul_result_o[7] = imul_result_o_7_sv2v_reg;
  assign imul_result_o[6] = imul_result_o_6_sv2v_reg;
  assign imul_result_o[5] = imul_result_o_5_sv2v_reg;
  assign imul_result_o[4] = imul_result_o_4_sv2v_reg;
  assign imul_result_o[3] = imul_result_o_3_sv2v_reg;
  assign imul_result_o[2] = imul_result_o_2_sv2v_reg;
  assign imul_result_o[1] = imul_result_o_1_sv2v_reg;
  assign imul_result_o[0] = imul_result_o_0_sv2v_reg;
  assign fma1_v_o = fma1_v_o_sv2v_reg;
  assign fma1_rm_o[2] = fma1_rm_o_2_sv2v_reg;
  assign fma1_rm_o[1] = fma1_rm_o_1_sv2v_reg;
  assign fma1_rm_o[0] = fma1_rm_o_0_sv2v_reg;
  assign imul_v_o = imul_v_o_sv2v_reg;
  assign out_sig_o[26] = out_sig_o_26_sv2v_reg;
  assign out_sig_o[25] = out_sig_o_25_sv2v_reg;
  assign out_sig_o[24] = out_sig_o_24_sv2v_reg;
  assign out_sig_o[23] = out_sig_o_23_sv2v_reg;
  assign out_sig_o[22] = out_sig_o_22_sv2v_reg;
  assign out_sig_o[21] = out_sig_o_21_sv2v_reg;
  assign out_sig_o[20] = out_sig_o_20_sv2v_reg;
  assign out_sig_o[19] = out_sig_o_19_sv2v_reg;
  assign out_sig_o[18] = out_sig_o_18_sv2v_reg;
  assign out_sig_o[17] = out_sig_o_17_sv2v_reg;
  assign out_sig_o[16] = out_sig_o_16_sv2v_reg;
  assign out_sig_o[15] = out_sig_o_15_sv2v_reg;
  assign out_sig_o[14] = out_sig_o_14_sv2v_reg;
  assign out_sig_o[13] = out_sig_o_13_sv2v_reg;
  assign out_sig_o[12] = out_sig_o_12_sv2v_reg;
  assign out_sig_o[11] = out_sig_o_11_sv2v_reg;
  assign out_sig_o[10] = out_sig_o_10_sv2v_reg;
  assign out_sig_o[9] = out_sig_o_9_sv2v_reg;
  assign out_sig_o[8] = out_sig_o_8_sv2v_reg;
  assign out_sig_o[7] = out_sig_o_7_sv2v_reg;
  assign out_sig_o[6] = out_sig_o_6_sv2v_reg;
  assign out_sig_o[5] = out_sig_o_5_sv2v_reg;
  assign out_sig_o[4] = out_sig_o_4_sv2v_reg;
  assign out_sig_o[3] = out_sig_o_3_sv2v_reg;
  assign out_sig_o[2] = out_sig_o_2_sv2v_reg;
  assign out_sig_o[1] = out_sig_o_1_sv2v_reg;
  assign out_sig_o[0] = out_sig_o_0_sv2v_reg;
  assign invalidExc_o = invalidExc_o_sv2v_reg;
  assign out_isNaN_o = out_isNaN_o_sv2v_reg;
  assign out_isInf_o = out_isInf_o_sv2v_reg;
  assign out_isZero_o = out_isZero_o_sv2v_reg;
  assign out_sign_o = out_sign_o_sv2v_reg;
  assign out_sExp_o[9] = out_sExp_o_9_sv2v_reg;
  assign out_sExp_o[8] = out_sExp_o_8_sv2v_reg;
  assign out_sExp_o[7] = out_sExp_o_7_sv2v_reg;
  assign out_sExp_o[6] = out_sExp_o_6_sv2v_reg;
  assign out_sExp_o[5] = out_sExp_o_5_sv2v_reg;
  assign out_sExp_o[4] = out_sExp_o_4_sv2v_reg;
  assign out_sExp_o[3] = out_sExp_o_3_sv2v_reg;
  assign out_sExp_o[2] = out_sExp_o_2_sv2v_reg;
  assign out_sExp_o[1] = out_sExp_o_1_sv2v_reg;
  assign out_sExp_o[0] = out_sExp_o_0_sv2v_reg;
  assign N18 = N14 & N15;
  assign N19 = N16 & N17;
  assign N20 = N18 & N19;
  assign N21 = fpu_float_op_i[3] | fpu_float_op_i[2];
  assign N22 = fpu_float_op_i[1] | N17;
  assign N23 = N21 | N22;
  assign N25 = N16 | fpu_float_op_i[0];
  assign N26 = N21 | N25;
  assign N28 = N14 | fpu_float_op_i[2];
  assign N29 = N16 | N17;
  assign N30 = N28 | N29;
  assign N32 = N14 | N15;
  assign N33 = fpu_float_op_i[1] | fpu_float_op_i[0];
  assign N34 = N32 | N33;
  assign N36 = N32 | N22;
  assign N38 = N32 | N25;
  assign N40 = N14 & fpu_float_op_i[1];
  assign N41 = N40 & fpu_float_op_i[0];
  assign N42 = fpu_float_op_i[2] & fpu_float_op_i[1];
  assign N43 = N42 & fpu_float_op_i[0];
  assign N44 = fpu_float_op_i[3] & N15;
  assign N45 = N44 & N16;
  assign N46 = N14 & fpu_float_op_i[2];
  assign N47 = N44 & N17;

  mulAddRecFNToRaw_expWidth8_sigWidth24
  mulAdd0
  (
    .control(1'b1),
    .op(fma_op_li),
    .a(fma_a_li),
    .b(fma_b_li),
    .c(fma_c_li),
    .roundingMode(fp_rm_i),
    .invalidExc(invalidExc),
    .out_isNaN(out_isNaN),
    .out_isInf(out_isInf),
    .out_isZero(out_isZero),
    .out_sign(out_sign),
    .out_sExp(out_sExp),
    .out_sig(out_sig),
    .out_imul(out_imul)
  );

  assign { N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49 } = (N0)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                   (N1)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                   (N3)? fp_rs2_i : 
                                                                                                                                                                                   (N4)? fp_rs2_i : 
                                                                                                                                                                                   (N5)? fp_rs2_i : 
                                                                                                                                                                                   (N6)? fp_rs2_i : 
                                                                                                                                                                                   (N7)? fp_rs2_i : 
                                                                                                                                                                                   (N8)? fp_rs2_i : 1'b0;
  assign N0 = N20;
  assign N1 = N24;
  assign N3 = N27;
  assign N4 = N31;
  assign N5 = N35;
  assign N6 = N37;
  assign N7 = N39;
  assign N8 = N48;
  assign { N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82 } = (N0)? fp_rs2_i : 
                                                                                                                                                                                                  (N1)? fp_rs2_i : 
                                                                                                                                                                                                  (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                  (N4)? fp_rs3_i : 
                                                                                                                                                                                                  (N5)? fp_rs3_i : 
                                                                                                                                                                                                  (N6)? fp_rs3_i : 
                                                                                                                                                                                                  (N7)? fp_rs3_i : 
                                                                                                                                                                                                  (N8)? fp_rs3_i : 1'b0;
  assign { N116, N115 } = (N0)? { 1'b0, 1'b0 } : 
                          (N1)? { 1'b0, 1'b1 } : 
                          (N3)? { 1'b0, 1'b0 } : 
                          (N4)? { 1'b0, 1'b0 } : 
                          (N5)? { 1'b0, 1'b1 } : 
                          (N6)? { 1'b1, 1'b0 } : 
                          (N7)? { 1'b1, 1'b1 } : 
                          (N8)? { 1'b0, 1'b0 } : 1'b0;
  assign N117 = (N0)? 1'b1 : 
                (N1)? 1'b1 : 
                (N3)? 1'b1 : 
                (N4)? 1'b1 : 
                (N5)? 1'b1 : 
                (N6)? 1'b1 : 
                (N7)? 1'b1 : 
                (N8)? 1'b0 : 1'b0;
  assign fma_a_li = (N9)? { 1'b0, imul_rs1_i } : 
                    (N10)? fp_rs1_i : 1'b0;
  assign N9 = fma_op_li[2];
  assign N10 = N123;
  assign fma_b_li = (N9)? { 1'b0, imul_rs2_i } : 
                    (N10)? { N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49 } : 1'b0;
  assign fma_c_li = (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                    (N10)? { N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82 } : 1'b0;
  assign fma_op_li[1:0] = (N9)? { 1'b0, 1'b0 } : 
                          (N10)? { N116, N115 } : 1'b0;
  assign is_fma_op = (N9)? 1'b0 : 
                     (N10)? N117 : 1'b0;
  assign N124 = (N11)? 1'b1 : 
                (N12)? 1'b0 : 1'b0;
  assign N11 = N118;
  assign N12 = stall_fpu1_i;
  assign N125 = (N11)? N122 : 
                (N12)? 1'b0 : 1'b0;
  assign N126 = (N13)? 1'b0 : 
                (N129)? N122 : 
                (N120)? 1'b0 : 1'b0;
  assign N13 = reset_i;
  assign N127 = (N13)? 1'b0 : 
                (N129)? imul_v_i : 
                (N120)? 1'b0 : 1'b0;
  assign fma_op_li[2] = imul_v_i;
  assign N14 = ~fpu_float_op_i[3];
  assign N15 = ~fpu_float_op_i[2];
  assign N16 = ~fpu_float_op_i[1];
  assign N17 = ~fpu_float_op_i[0];
  assign N24 = ~N23;
  assign N27 = ~N26;
  assign N31 = ~N30;
  assign N35 = ~N34;
  assign N37 = ~N36;
  assign N39 = ~N38;
  assign N48 = N41 | N132;
  assign N132 = N43 | N131;
  assign N131 = N45 | N130;
  assign N130 = N46 | N47;
  assign N118 = ~stall_fpu1_i;
  assign N119 = N118 | reset_i;
  assign N120 = ~N119;
  assign N121 = fp_v_i & is_fma_op;
  assign N122 = fp_v_i & is_fma_op;
  assign N123 = ~imul_v_i;
  assign N128 = ~reset_i;
  assign N129 = N118 & N128;

  always @(posedge clk_i) begin
    if(N127) begin
      imul_result_o_31_sv2v_reg <= out_imul[31];
      imul_result_o_30_sv2v_reg <= out_imul[30];
      imul_result_o_29_sv2v_reg <= out_imul[29];
      imul_result_o_28_sv2v_reg <= out_imul[28];
      imul_result_o_27_sv2v_reg <= out_imul[27];
      imul_result_o_26_sv2v_reg <= out_imul[26];
      imul_result_o_25_sv2v_reg <= out_imul[25];
      imul_result_o_24_sv2v_reg <= out_imul[24];
      imul_result_o_23_sv2v_reg <= out_imul[23];
      imul_result_o_22_sv2v_reg <= out_imul[22];
      imul_result_o_21_sv2v_reg <= out_imul[21];
      imul_result_o_20_sv2v_reg <= out_imul[20];
      imul_result_o_19_sv2v_reg <= out_imul[19];
      imul_result_o_18_sv2v_reg <= out_imul[18];
      imul_result_o_17_sv2v_reg <= out_imul[17];
      imul_result_o_16_sv2v_reg <= out_imul[16];
      imul_result_o_15_sv2v_reg <= out_imul[15];
      imul_result_o_14_sv2v_reg <= out_imul[14];
      imul_result_o_13_sv2v_reg <= out_imul[13];
      imul_result_o_12_sv2v_reg <= out_imul[12];
      imul_result_o_11_sv2v_reg <= out_imul[11];
      imul_result_o_10_sv2v_reg <= out_imul[10];
      imul_result_o_9_sv2v_reg <= out_imul[9];
      imul_result_o_8_sv2v_reg <= out_imul[8];
      imul_result_o_7_sv2v_reg <= out_imul[7];
      imul_result_o_6_sv2v_reg <= out_imul[6];
      imul_result_o_5_sv2v_reg <= out_imul[5];
      imul_result_o_4_sv2v_reg <= out_imul[4];
      imul_result_o_3_sv2v_reg <= out_imul[3];
      imul_result_o_2_sv2v_reg <= out_imul[2];
      imul_result_o_1_sv2v_reg <= out_imul[1];
      imul_result_o_0_sv2v_reg <= out_imul[0];
    end 
    if(reset_i) begin
      fma1_v_o_sv2v_reg <= 1'b0;
      imul_v_o_sv2v_reg <= 1'b0;
    end else if(N124) begin
      fma1_v_o_sv2v_reg <= N121;
      imul_v_o_sv2v_reg <= imul_v_i;
    end 
    if(reset_i) begin
      fma1_rm_o_2_sv2v_reg <= 1'b1;
      fma1_rm_o_1_sv2v_reg <= 1'b1;
      fma1_rm_o_0_sv2v_reg <= 1'b1;
    end else if(N125) begin
      fma1_rm_o_2_sv2v_reg <= fp_rm_i[2];
      fma1_rm_o_1_sv2v_reg <= fp_rm_i[1];
      fma1_rm_o_0_sv2v_reg <= fp_rm_i[0];
    end 
    if(N126) begin
      out_sig_o_26_sv2v_reg <= out_sig[26];
      out_sig_o_25_sv2v_reg <= out_sig[25];
      out_sig_o_24_sv2v_reg <= out_sig[24];
      out_sig_o_23_sv2v_reg <= out_sig[23];
      out_sig_o_22_sv2v_reg <= out_sig[22];
      out_sig_o_21_sv2v_reg <= out_sig[21];
      out_sig_o_20_sv2v_reg <= out_sig[20];
      out_sig_o_19_sv2v_reg <= out_sig[19];
      out_sig_o_18_sv2v_reg <= out_sig[18];
      out_sig_o_17_sv2v_reg <= out_sig[17];
      out_sig_o_16_sv2v_reg <= out_sig[16];
      out_sig_o_15_sv2v_reg <= out_sig[15];
      out_sig_o_14_sv2v_reg <= out_sig[14];
      out_sig_o_13_sv2v_reg <= out_sig[13];
      out_sig_o_12_sv2v_reg <= out_sig[12];
      out_sig_o_11_sv2v_reg <= out_sig[11];
      out_sig_o_10_sv2v_reg <= out_sig[10];
      out_sig_o_9_sv2v_reg <= out_sig[9];
      out_sig_o_8_sv2v_reg <= out_sig[8];
      out_sig_o_7_sv2v_reg <= out_sig[7];
      out_sig_o_6_sv2v_reg <= out_sig[6];
      out_sig_o_5_sv2v_reg <= out_sig[5];
      out_sig_o_4_sv2v_reg <= out_sig[4];
      out_sig_o_3_sv2v_reg <= out_sig[3];
      out_sig_o_2_sv2v_reg <= out_sig[2];
      out_sig_o_1_sv2v_reg <= out_sig[1];
      out_sig_o_0_sv2v_reg <= out_sig[0];
      invalidExc_o_sv2v_reg <= invalidExc;
      out_isNaN_o_sv2v_reg <= out_isNaN;
      out_isInf_o_sv2v_reg <= out_isInf;
      out_isZero_o_sv2v_reg <= out_isZero;
      out_sign_o_sv2v_reg <= out_sign;
      out_sExp_o_9_sv2v_reg <= out_sExp[9];
      out_sExp_o_8_sv2v_reg <= out_sExp[8];
      out_sExp_o_7_sv2v_reg <= out_sExp[7];
      out_sExp_o_6_sv2v_reg <= out_sExp[6];
      out_sExp_o_5_sv2v_reg <= out_sExp[5];
      out_sExp_o_4_sv2v_reg <= out_sExp[4];
      out_sExp_o_3_sv2v_reg <= out_sExp[3];
      out_sExp_o_2_sv2v_reg <= out_sExp[2];
      out_sExp_o_1_sv2v_reg <= out_sExp[1];
      out_sExp_o_0_sv2v_reg <= out_sExp[0];
    end 
  end


endmodule



module reverse_width25
(
  in,
  out
);

  input [24:0] in;
  output [24:0] out;
  wire [24:0] out;
  assign out[24] = in[0];
  assign out[23] = in[1];
  assign out[22] = in[2];
  assign out[21] = in[3];
  assign out[20] = in[4];
  assign out[19] = in[5];
  assign out[18] = in[6];
  assign out[17] = in[7];
  assign out[16] = in[8];
  assign out[15] = in[9];
  assign out[14] = in[10];
  assign out[13] = in[11];
  assign out[12] = in[12];
  assign out[11] = in[13];
  assign out[10] = in[14];
  assign out[9] = in[15];
  assign out[8] = in[16];
  assign out[7] = in[17];
  assign out[6] = in[18];
  assign out[5] = in[19];
  assign out[4] = in[20];
  assign out[3] = in[21];
  assign out[2] = in[22];
  assign out[1] = in[23];
  assign out[0] = in[24];

endmodule



module lowMaskLoHi_inWidth9_topBound105_bottomBound130
(
  in,
  out
);

  input [8:0] in;
  output [24:0] out;
  wire [24:0] out,reverseOut;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,
  sv2v_dc_6,sv2v_dc_7,sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,
  sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,
  sv2v_dc_21,sv2v_dc_22,sv2v_dc_23,sv2v_dc_24,sv2v_dc_25,sv2v_dc_26,sv2v_dc_27,
  sv2v_dc_28,sv2v_dc_29,sv2v_dc_30,sv2v_dc_31,sv2v_dc_32,sv2v_dc_33,sv2v_dc_34,
  sv2v_dc_35,sv2v_dc_36,sv2v_dc_37,sv2v_dc_38,sv2v_dc_39,sv2v_dc_40,sv2v_dc_41,sv2v_dc_42,
  sv2v_dc_43,sv2v_dc_44,sv2v_dc_45,sv2v_dc_46,sv2v_dc_47,sv2v_dc_48,sv2v_dc_49,
  sv2v_dc_50,sv2v_dc_51,sv2v_dc_52,sv2v_dc_53,sv2v_dc_54,sv2v_dc_55,sv2v_dc_56,
  sv2v_dc_57,sv2v_dc_58,sv2v_dc_59,sv2v_dc_60,sv2v_dc_61,sv2v_dc_62,sv2v_dc_63,
  sv2v_dc_64,sv2v_dc_65,sv2v_dc_66,sv2v_dc_67,sv2v_dc_68,sv2v_dc_69,sv2v_dc_70,sv2v_dc_71,
  sv2v_dc_72,sv2v_dc_73,sv2v_dc_74,sv2v_dc_75,sv2v_dc_76,sv2v_dc_77,sv2v_dc_78,
  sv2v_dc_79,sv2v_dc_80,sv2v_dc_81,sv2v_dc_82,sv2v_dc_83,sv2v_dc_84,sv2v_dc_85,
  sv2v_dc_86,sv2v_dc_87,sv2v_dc_88,sv2v_dc_89,sv2v_dc_90,sv2v_dc_91,sv2v_dc_92,
  sv2v_dc_93,sv2v_dc_94,sv2v_dc_95,sv2v_dc_96,sv2v_dc_97,sv2v_dc_98,sv2v_dc_99,sv2v_dc_100,
  sv2v_dc_101,sv2v_dc_102,sv2v_dc_103,sv2v_dc_104,sv2v_dc_105,sv2v_dc_106,
  sv2v_dc_107,sv2v_dc_108,sv2v_dc_109,sv2v_dc_110,sv2v_dc_111,sv2v_dc_112,sv2v_dc_113,
  sv2v_dc_114,sv2v_dc_115,sv2v_dc_116,sv2v_dc_117,sv2v_dc_118,sv2v_dc_119,sv2v_dc_120,
  sv2v_dc_121,sv2v_dc_122,sv2v_dc_123,sv2v_dc_124,sv2v_dc_125,sv2v_dc_126,
  sv2v_dc_127,sv2v_dc_128,sv2v_dc_129,sv2v_dc_130,sv2v_dc_131,sv2v_dc_132,sv2v_dc_133,
  sv2v_dc_134,sv2v_dc_135,sv2v_dc_136,sv2v_dc_137,sv2v_dc_138,sv2v_dc_139,sv2v_dc_140,
  sv2v_dc_141,sv2v_dc_142,sv2v_dc_143,sv2v_dc_144,sv2v_dc_145,sv2v_dc_146,
  sv2v_dc_147,sv2v_dc_148,sv2v_dc_149,sv2v_dc_150,sv2v_dc_151,sv2v_dc_152,sv2v_dc_153,
  sv2v_dc_154,sv2v_dc_155,sv2v_dc_156,sv2v_dc_157,sv2v_dc_158,sv2v_dc_159,sv2v_dc_160,
  sv2v_dc_161,sv2v_dc_162,sv2v_dc_163,sv2v_dc_164,sv2v_dc_165,sv2v_dc_166,
  sv2v_dc_167,sv2v_dc_168,sv2v_dc_169,sv2v_dc_170,sv2v_dc_171,sv2v_dc_172,sv2v_dc_173,
  sv2v_dc_174,sv2v_dc_175,sv2v_dc_176,sv2v_dc_177,sv2v_dc_178,sv2v_dc_179,sv2v_dc_180,
  sv2v_dc_181,sv2v_dc_182,sv2v_dc_183,sv2v_dc_184,sv2v_dc_185,sv2v_dc_186,
  sv2v_dc_187,sv2v_dc_188,sv2v_dc_189,sv2v_dc_190,sv2v_dc_191,sv2v_dc_192,sv2v_dc_193,
  sv2v_dc_194,sv2v_dc_195,sv2v_dc_196,sv2v_dc_197,sv2v_dc_198,sv2v_dc_199,sv2v_dc_200,
  sv2v_dc_201,sv2v_dc_202,sv2v_dc_203,sv2v_dc_204,sv2v_dc_205,sv2v_dc_206,
  sv2v_dc_207,sv2v_dc_208,sv2v_dc_209,sv2v_dc_210,sv2v_dc_211,sv2v_dc_212,sv2v_dc_213,
  sv2v_dc_214,sv2v_dc_215,sv2v_dc_216,sv2v_dc_217,sv2v_dc_218,sv2v_dc_219,sv2v_dc_220,
  sv2v_dc_221,sv2v_dc_222,sv2v_dc_223,sv2v_dc_224,sv2v_dc_225,sv2v_dc_226,
  sv2v_dc_227,sv2v_dc_228,sv2v_dc_229,sv2v_dc_230,sv2v_dc_231,sv2v_dc_232,sv2v_dc_233,
  sv2v_dc_234,sv2v_dc_235,sv2v_dc_236,sv2v_dc_237,sv2v_dc_238,sv2v_dc_239,sv2v_dc_240,
  sv2v_dc_241,sv2v_dc_242,sv2v_dc_243,sv2v_dc_244,sv2v_dc_245,sv2v_dc_246,
  sv2v_dc_247,sv2v_dc_248,sv2v_dc_249,sv2v_dc_250,sv2v_dc_251,sv2v_dc_252,sv2v_dc_253,
  sv2v_dc_254,sv2v_dc_255,sv2v_dc_256,sv2v_dc_257,sv2v_dc_258,sv2v_dc_259,sv2v_dc_260,
  sv2v_dc_261,sv2v_dc_262,sv2v_dc_263,sv2v_dc_264,sv2v_dc_265,sv2v_dc_266,
  sv2v_dc_267,sv2v_dc_268,sv2v_dc_269,sv2v_dc_270,sv2v_dc_271,sv2v_dc_272,sv2v_dc_273,
  sv2v_dc_274,sv2v_dc_275,sv2v_dc_276,sv2v_dc_277,sv2v_dc_278,sv2v_dc_279,sv2v_dc_280,
  sv2v_dc_281,sv2v_dc_282,sv2v_dc_283,sv2v_dc_284,sv2v_dc_285,sv2v_dc_286,
  sv2v_dc_287,sv2v_dc_288,sv2v_dc_289,sv2v_dc_290,sv2v_dc_291,sv2v_dc_292,sv2v_dc_293,
  sv2v_dc_294,sv2v_dc_295,sv2v_dc_296,sv2v_dc_297,sv2v_dc_298,sv2v_dc_299,sv2v_dc_300,
  sv2v_dc_301,sv2v_dc_302,sv2v_dc_303,sv2v_dc_304,sv2v_dc_305,sv2v_dc_306,
  sv2v_dc_307,sv2v_dc_308,sv2v_dc_309,sv2v_dc_310,sv2v_dc_311,sv2v_dc_312,sv2v_dc_313,
  sv2v_dc_314,sv2v_dc_315,sv2v_dc_316,sv2v_dc_317,sv2v_dc_318,sv2v_dc_319,sv2v_dc_320,
  sv2v_dc_321,sv2v_dc_322,sv2v_dc_323,sv2v_dc_324,sv2v_dc_325,sv2v_dc_326,
  sv2v_dc_327,sv2v_dc_328,sv2v_dc_329,sv2v_dc_330,sv2v_dc_331,sv2v_dc_332,sv2v_dc_333,
  sv2v_dc_334,sv2v_dc_335,sv2v_dc_336,sv2v_dc_337,sv2v_dc_338,sv2v_dc_339,sv2v_dc_340,
  sv2v_dc_341,sv2v_dc_342,sv2v_dc_343,sv2v_dc_344,sv2v_dc_345,sv2v_dc_346,
  sv2v_dc_347,sv2v_dc_348,sv2v_dc_349,sv2v_dc_350,sv2v_dc_351,sv2v_dc_352,sv2v_dc_353,
  sv2v_dc_354,sv2v_dc_355,sv2v_dc_356,sv2v_dc_357,sv2v_dc_358,sv2v_dc_359,sv2v_dc_360,
  sv2v_dc_361,sv2v_dc_362,sv2v_dc_363,sv2v_dc_364,sv2v_dc_365,sv2v_dc_366,
  sv2v_dc_367,sv2v_dc_368,sv2v_dc_369,sv2v_dc_370,sv2v_dc_371,sv2v_dc_372,sv2v_dc_373,
  sv2v_dc_374,sv2v_dc_375,sv2v_dc_376,sv2v_dc_377,sv2v_dc_378,sv2v_dc_379,sv2v_dc_380,
  sv2v_dc_381,sv2v_dc_382;

  reverse_width25
  reverse
  (
    .in(reverseOut),
    .out(out)
  );

  assign { sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25, sv2v_dc_26, sv2v_dc_27, sv2v_dc_28, sv2v_dc_29, sv2v_dc_30, sv2v_dc_31, sv2v_dc_32, sv2v_dc_33, sv2v_dc_34, sv2v_dc_35, sv2v_dc_36, sv2v_dc_37, sv2v_dc_38, sv2v_dc_39, sv2v_dc_40, sv2v_dc_41, sv2v_dc_42, sv2v_dc_43, sv2v_dc_44, sv2v_dc_45, sv2v_dc_46, sv2v_dc_47, sv2v_dc_48, sv2v_dc_49, sv2v_dc_50, sv2v_dc_51, sv2v_dc_52, sv2v_dc_53, sv2v_dc_54, sv2v_dc_55, sv2v_dc_56, sv2v_dc_57, sv2v_dc_58, sv2v_dc_59, sv2v_dc_60, sv2v_dc_61, sv2v_dc_62, sv2v_dc_63, sv2v_dc_64, sv2v_dc_65, sv2v_dc_66, sv2v_dc_67, sv2v_dc_68, sv2v_dc_69, sv2v_dc_70, sv2v_dc_71, sv2v_dc_72, sv2v_dc_73, sv2v_dc_74, sv2v_dc_75, sv2v_dc_76, sv2v_dc_77, sv2v_dc_78, sv2v_dc_79, sv2v_dc_80, sv2v_dc_81, sv2v_dc_82, sv2v_dc_83, sv2v_dc_84, sv2v_dc_85, sv2v_dc_86, sv2v_dc_87, sv2v_dc_88, sv2v_dc_89, sv2v_dc_90, sv2v_dc_91, sv2v_dc_92, sv2v_dc_93, sv2v_dc_94, sv2v_dc_95, sv2v_dc_96, sv2v_dc_97, sv2v_dc_98, sv2v_dc_99, sv2v_dc_100, sv2v_dc_101, sv2v_dc_102, sv2v_dc_103, sv2v_dc_104, sv2v_dc_105, sv2v_dc_106, sv2v_dc_107, sv2v_dc_108, sv2v_dc_109, sv2v_dc_110, sv2v_dc_111, sv2v_dc_112, sv2v_dc_113, sv2v_dc_114, sv2v_dc_115, sv2v_dc_116, sv2v_dc_117, sv2v_dc_118, sv2v_dc_119, sv2v_dc_120, sv2v_dc_121, sv2v_dc_122, sv2v_dc_123, sv2v_dc_124, sv2v_dc_125, sv2v_dc_126, sv2v_dc_127, sv2v_dc_128, sv2v_dc_129, sv2v_dc_130, sv2v_dc_131, sv2v_dc_132, sv2v_dc_133, sv2v_dc_134, sv2v_dc_135, sv2v_dc_136, sv2v_dc_137, sv2v_dc_138, sv2v_dc_139, sv2v_dc_140, sv2v_dc_141, sv2v_dc_142, sv2v_dc_143, sv2v_dc_144, sv2v_dc_145, sv2v_dc_146, sv2v_dc_147, sv2v_dc_148, sv2v_dc_149, sv2v_dc_150, sv2v_dc_151, sv2v_dc_152, sv2v_dc_153, sv2v_dc_154, sv2v_dc_155, sv2v_dc_156, sv2v_dc_157, sv2v_dc_158, sv2v_dc_159, sv2v_dc_160, sv2v_dc_161, sv2v_dc_162, sv2v_dc_163, sv2v_dc_164, sv2v_dc_165, sv2v_dc_166, sv2v_dc_167, sv2v_dc_168, sv2v_dc_169, sv2v_dc_170, sv2v_dc_171, sv2v_dc_172, sv2v_dc_173, sv2v_dc_174, sv2v_dc_175, sv2v_dc_176, sv2v_dc_177, sv2v_dc_178, sv2v_dc_179, sv2v_dc_180, sv2v_dc_181, sv2v_dc_182, sv2v_dc_183, sv2v_dc_184, sv2v_dc_185, sv2v_dc_186, sv2v_dc_187, sv2v_dc_188, sv2v_dc_189, sv2v_dc_190, sv2v_dc_191, sv2v_dc_192, sv2v_dc_193, sv2v_dc_194, sv2v_dc_195, sv2v_dc_196, sv2v_dc_197, sv2v_dc_198, sv2v_dc_199, sv2v_dc_200, sv2v_dc_201, sv2v_dc_202, sv2v_dc_203, sv2v_dc_204, sv2v_dc_205, sv2v_dc_206, sv2v_dc_207, sv2v_dc_208, sv2v_dc_209, sv2v_dc_210, sv2v_dc_211, sv2v_dc_212, sv2v_dc_213, sv2v_dc_214, sv2v_dc_215, sv2v_dc_216, sv2v_dc_217, sv2v_dc_218, sv2v_dc_219, sv2v_dc_220, sv2v_dc_221, sv2v_dc_222, sv2v_dc_223, sv2v_dc_224, sv2v_dc_225, sv2v_dc_226, sv2v_dc_227, sv2v_dc_228, sv2v_dc_229, sv2v_dc_230, sv2v_dc_231, sv2v_dc_232, sv2v_dc_233, sv2v_dc_234, sv2v_dc_235, sv2v_dc_236, sv2v_dc_237, sv2v_dc_238, sv2v_dc_239, sv2v_dc_240, sv2v_dc_241, sv2v_dc_242, sv2v_dc_243, sv2v_dc_244, sv2v_dc_245, sv2v_dc_246, sv2v_dc_247, sv2v_dc_248, sv2v_dc_249, sv2v_dc_250, sv2v_dc_251, sv2v_dc_252, sv2v_dc_253, sv2v_dc_254, sv2v_dc_255, sv2v_dc_256, sv2v_dc_257, sv2v_dc_258, sv2v_dc_259, sv2v_dc_260, sv2v_dc_261, sv2v_dc_262, sv2v_dc_263, sv2v_dc_264, sv2v_dc_265, sv2v_dc_266, sv2v_dc_267, sv2v_dc_268, sv2v_dc_269, sv2v_dc_270, sv2v_dc_271, sv2v_dc_272, sv2v_dc_273, sv2v_dc_274, sv2v_dc_275, sv2v_dc_276, sv2v_dc_277, sv2v_dc_278, sv2v_dc_279, sv2v_dc_280, sv2v_dc_281, sv2v_dc_282, sv2v_dc_283, sv2v_dc_284, sv2v_dc_285, sv2v_dc_286, sv2v_dc_287, sv2v_dc_288, sv2v_dc_289, sv2v_dc_290, sv2v_dc_291, sv2v_dc_292, sv2v_dc_293, sv2v_dc_294, sv2v_dc_295, sv2v_dc_296, sv2v_dc_297, sv2v_dc_298, sv2v_dc_299, sv2v_dc_300, sv2v_dc_301, sv2v_dc_302, sv2v_dc_303, sv2v_dc_304, sv2v_dc_305, sv2v_dc_306, sv2v_dc_307, sv2v_dc_308, sv2v_dc_309, sv2v_dc_310, sv2v_dc_311, sv2v_dc_312, sv2v_dc_313, sv2v_dc_314, sv2v_dc_315, sv2v_dc_316, sv2v_dc_317, sv2v_dc_318, sv2v_dc_319, sv2v_dc_320, sv2v_dc_321, sv2v_dc_322, sv2v_dc_323, sv2v_dc_324, sv2v_dc_325, sv2v_dc_326, sv2v_dc_327, sv2v_dc_328, sv2v_dc_329, sv2v_dc_330, sv2v_dc_331, sv2v_dc_332, sv2v_dc_333, sv2v_dc_334, sv2v_dc_335, sv2v_dc_336, sv2v_dc_337, sv2v_dc_338, sv2v_dc_339, sv2v_dc_340, sv2v_dc_341, sv2v_dc_342, sv2v_dc_343, sv2v_dc_344, sv2v_dc_345, sv2v_dc_346, sv2v_dc_347, sv2v_dc_348, sv2v_dc_349, sv2v_dc_350, sv2v_dc_351, sv2v_dc_352, sv2v_dc_353, sv2v_dc_354, sv2v_dc_355, sv2v_dc_356, sv2v_dc_357, sv2v_dc_358, sv2v_dc_359, sv2v_dc_360, sv2v_dc_361, sv2v_dc_362, sv2v_dc_363, sv2v_dc_364, sv2v_dc_365, sv2v_dc_366, sv2v_dc_367, sv2v_dc_368, sv2v_dc_369, sv2v_dc_370, sv2v_dc_371, sv2v_dc_372, sv2v_dc_373, sv2v_dc_374, sv2v_dc_375, sv2v_dc_376, sv2v_dc_377, sv2v_dc_378, sv2v_dc_379, sv2v_dc_380, sv2v_dc_381, sv2v_dc_382, reverseOut } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { N0, N1, N2, N3, N4, N5, N6, N7, N8 };
  assign N0 = ~in[8];
  assign N1 = ~in[7];
  assign N2 = ~in[6];
  assign N3 = ~in[5];
  assign N4 = ~in[4];
  assign N5 = ~in[3];
  assign N6 = ~in[2];
  assign N7 = ~in[1];
  assign N8 = ~in[0];

endmodule



module roundAnyRawFNToRecFN_inExpWidth8_inSigWidth26_outExpWidth8_outSigWidth24_options0
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [9:0] in_sExp;
  input [26:0] in_sig;
  input [2:0] roundingMode;
  output [32:0] out;
  output [4:0] exceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [32:0] out;
  wire [4:0] exceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,exceptionFlags_4_,
  exceptionFlags_3_,roundMagUp,isNaNOut,_0_net__8_,\genblk2.roundPosBit ,\genblk2.anyRoundExtra ,
  \genblk2.anyRound ,\genblk2.roundIncr ,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,
  N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,
  N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,common_overflow,common_totalUnderflow,
  \genblk2.unboundedRange_roundPosBit ,\genblk2.unboundedRange_anyRound ,
  \genblk2.unboundedRange_roundIncr ,\genblk2.roundCarry ,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  common_underflow,common_inexact,notNaN_isSpecialInfOut,commonCase,
  overflow_roundMagUp,pegMinNonzeroMagOut,pegMaxFiniteMagOut,notNaN_isInfOut,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465;
  wire [24:0] \genblk2.genblk1.roundMask_main ;
  wire [2:2] \genblk2.roundMask ;
  wire [26:0] \genblk2.roundPosMask ;
  wire [25:0] \genblk2.roundedSig ;
  wire [10:0] \genblk2.sRoundedExp ;
  wire [22:0] common_fractOut;
  assign exceptionFlags_4_ = invalidExc;
  assign exceptionFlags[4] = exceptionFlags_4_;
  assign exceptionFlags_3_ = infiniteExc;
  assign exceptionFlags[3] = exceptionFlags_3_;

  lowMaskLoHi_inWidth9_topBound105_bottomBound130
  \genblk2.genblk1.lowMask_roundMask 
  (
    .in({ _0_net__8_, in_sExp[7:0] }),
    .out(\genblk2.genblk1.roundMask_main )
  );

  assign common_overflow = $signed(\genblk2.sRoundedExp [10:7]) >= $signed({ 1'b0, 1'b1, 1'b1 });
  assign common_totalUnderflow = $signed(\genblk2.sRoundedExp ) < $signed({ 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 });
  assign N174 = $signed(in_sExp[9:8]) <= $signed(1'b0);
  assign N210 = ~roundingMode[2];
  assign N211 = ~roundingMode[1];
  assign N212 = N211 | N210;
  assign N213 = roundingMode[0] | N212;
  assign N214 = ~N213;
  assign N215 = roundingMode[1] | N210;
  assign N216 = roundingMode[0] | N215;
  assign N217 = ~N216;
  assign N218 = roundingMode[1] | roundingMode[2];
  assign N219 = roundingMode[0] | N218;
  assign N220 = ~N219;
  assign N221 = N211 | roundingMode[2];
  assign N222 = roundingMode[0] | N221;
  assign N223 = ~N222;
  assign N224 = ~roundingMode[0];
  assign N225 = N224 | N221;
  assign N226 = ~N225;
  assign { N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67 } = { N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66 } + 1'b1;
  assign \genblk2.sRoundedExp  = { in_sExp[9:9], in_sExp } + \genblk2.roundedSig [25:24];
  assign { N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17 } = (N0)? { \genblk2.genblk1.roundMask_main [24:1], \genblk2.roundMask [2:2] } : 
                                                                                                                                           (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N15;
  assign { N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121 } = (N1)? \genblk2.roundPosMask [26:1] : 
                                                                                                                                                                          (N120)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = N119;
  assign \genblk2.roundedSig  = (N2)? { N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118 } : 
                                (N3)? { N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171 } : 1'b0;
  assign N2 = \genblk2.roundIncr ;
  assign N3 = N14;
  assign common_fractOut = (N4)? \genblk2.roundedSig [23:1] : 
                           (N5)? \genblk2.roundedSig [22:0] : 1'b0;
  assign N4 = in_sig[26];
  assign N5 = N172;
  assign \genblk2.unboundedRange_roundPosBit  = (N4)? in_sig[2] : 
                                                (N5)? in_sig[1] : 1'b0;
  assign \genblk2.roundCarry  = (N4)? \genblk2.roundedSig [25] : 
                                (N5)? \genblk2.roundedSig [24] : 1'b0;
  assign N173 = (N4)? \genblk2.genblk1.roundMask_main [1] : 
                (N5)? \genblk2.roundMask [2] : 1'b0;
  assign N177 = (N6)? N173 : 
                (N7)? 1'b0 : 1'b0;
  assign N6 = N175;
  assign N7 = N176;
  assign N178 = (N4)? \genblk2.genblk1.roundMask_main [2] : 
                (N5)? \genblk2.genblk1.roundMask_main [1] : 1'b0;
  assign N181 = (N8)? N180 : 
                (N9)? 1'b0 : 1'b0;
  assign N8 = control[0];
  assign N9 = N179;
  assign out[32] = (N10)? 1'b0 : 
                   (N11)? in_sign : 1'b0;
  assign N10 = isNaNOut;
  assign N11 = N431;
  assign N185 = (N12)? common_fractOut[22] : 
                (N184)? 1'b0 : 1'b0;
  assign N12 = N183;
  assign { N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188 } = (N13)? common_fractOut[21:0] : 
                                                                                                                                                  (N187)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N186;
  assign roundMagUp = N227 | N229;
  assign N227 = N223 & in_sign;
  assign N229 = N226 & N228;
  assign N228 = ~in_sign;
  assign isNaNOut = exceptionFlags_4_ | N231;
  assign N231 = N230 & in_isNaN;
  assign N230 = ~exceptionFlags_3_;
  assign _0_net__8_ = in_sExp[8] | 1'b0;
  assign \genblk2.roundMask [2] = \genblk2.genblk1.roundMask_main [0] | in_sig[26];
  assign \genblk2.roundPosMask [26] = N232 & \genblk2.genblk1.roundMask_main [24];
  assign N232 = ~1'b0;
  assign \genblk2.roundPosMask [25] = N233 & \genblk2.genblk1.roundMask_main [23];
  assign N233 = ~\genblk2.genblk1.roundMask_main [24];
  assign \genblk2.roundPosMask [24] = N234 & \genblk2.genblk1.roundMask_main [22];
  assign N234 = ~\genblk2.genblk1.roundMask_main [23];
  assign \genblk2.roundPosMask [23] = N235 & \genblk2.genblk1.roundMask_main [21];
  assign N235 = ~\genblk2.genblk1.roundMask_main [22];
  assign \genblk2.roundPosMask [22] = N236 & \genblk2.genblk1.roundMask_main [20];
  assign N236 = ~\genblk2.genblk1.roundMask_main [21];
  assign \genblk2.roundPosMask [21] = N237 & \genblk2.genblk1.roundMask_main [19];
  assign N237 = ~\genblk2.genblk1.roundMask_main [20];
  assign \genblk2.roundPosMask [20] = N238 & \genblk2.genblk1.roundMask_main [18];
  assign N238 = ~\genblk2.genblk1.roundMask_main [19];
  assign \genblk2.roundPosMask [19] = N239 & \genblk2.genblk1.roundMask_main [17];
  assign N239 = ~\genblk2.genblk1.roundMask_main [18];
  assign \genblk2.roundPosMask [18] = N240 & \genblk2.genblk1.roundMask_main [16];
  assign N240 = ~\genblk2.genblk1.roundMask_main [17];
  assign \genblk2.roundPosMask [17] = N241 & \genblk2.genblk1.roundMask_main [15];
  assign N241 = ~\genblk2.genblk1.roundMask_main [16];
  assign \genblk2.roundPosMask [16] = N242 & \genblk2.genblk1.roundMask_main [14];
  assign N242 = ~\genblk2.genblk1.roundMask_main [15];
  assign \genblk2.roundPosMask [15] = N243 & \genblk2.genblk1.roundMask_main [13];
  assign N243 = ~\genblk2.genblk1.roundMask_main [14];
  assign \genblk2.roundPosMask [14] = N244 & \genblk2.genblk1.roundMask_main [12];
  assign N244 = ~\genblk2.genblk1.roundMask_main [13];
  assign \genblk2.roundPosMask [13] = N245 & \genblk2.genblk1.roundMask_main [11];
  assign N245 = ~\genblk2.genblk1.roundMask_main [12];
  assign \genblk2.roundPosMask [12] = N246 & \genblk2.genblk1.roundMask_main [10];
  assign N246 = ~\genblk2.genblk1.roundMask_main [11];
  assign \genblk2.roundPosMask [11] = N247 & \genblk2.genblk1.roundMask_main [9];
  assign N247 = ~\genblk2.genblk1.roundMask_main [10];
  assign \genblk2.roundPosMask [10] = N248 & \genblk2.genblk1.roundMask_main [8];
  assign N248 = ~\genblk2.genblk1.roundMask_main [9];
  assign \genblk2.roundPosMask [9] = N249 & \genblk2.genblk1.roundMask_main [7];
  assign N249 = ~\genblk2.genblk1.roundMask_main [8];
  assign \genblk2.roundPosMask [8] = N250 & \genblk2.genblk1.roundMask_main [6];
  assign N250 = ~\genblk2.genblk1.roundMask_main [7];
  assign \genblk2.roundPosMask [7] = N251 & \genblk2.genblk1.roundMask_main [5];
  assign N251 = ~\genblk2.genblk1.roundMask_main [6];
  assign \genblk2.roundPosMask [6] = N252 & \genblk2.genblk1.roundMask_main [4];
  assign N252 = ~\genblk2.genblk1.roundMask_main [5];
  assign \genblk2.roundPosMask [5] = N253 & \genblk2.genblk1.roundMask_main [3];
  assign N253 = ~\genblk2.genblk1.roundMask_main [4];
  assign \genblk2.roundPosMask [4] = N254 & \genblk2.genblk1.roundMask_main [2];
  assign N254 = ~\genblk2.genblk1.roundMask_main [3];
  assign \genblk2.roundPosMask [3] = N255 & \genblk2.genblk1.roundMask_main [1];
  assign N255 = ~\genblk2.genblk1.roundMask_main [2];
  assign \genblk2.roundPosMask [2] = N256 & \genblk2.roundMask [2];
  assign N256 = ~\genblk2.genblk1.roundMask_main [1];
  assign \genblk2.roundPosMask [1] = N257 & 1'b1;
  assign N257 = ~\genblk2.roundMask [2];
  assign \genblk2.roundPosMask [0] = N258 & 1'b1;
  assign N258 = ~1'b1;
  assign \genblk2.roundPosBit  = N305 | N311;
  assign N305 = N303 | N304;
  assign N303 = N301 | N302;
  assign N301 = N299 | N300;
  assign N299 = N297 | N298;
  assign N297 = N295 | N296;
  assign N295 = N293 | N294;
  assign N293 = N291 | N292;
  assign N291 = N289 | N290;
  assign N289 = N287 | N288;
  assign N287 = N285 | N286;
  assign N285 = N283 | N284;
  assign N283 = N281 | N282;
  assign N281 = N279 | N280;
  assign N279 = N277 | N278;
  assign N277 = N275 | N276;
  assign N275 = N273 | N274;
  assign N273 = N271 | N272;
  assign N271 = N269 | N270;
  assign N269 = N267 | N268;
  assign N267 = N265 | N266;
  assign N265 = N263 | N264;
  assign N263 = N261 | N262;
  assign N261 = N259 | N260;
  assign N259 = in_sig[26] & \genblk2.roundPosMask [26];
  assign N260 = in_sig[25] & \genblk2.roundPosMask [25];
  assign N262 = in_sig[24] & \genblk2.roundPosMask [24];
  assign N264 = in_sig[23] & \genblk2.roundPosMask [23];
  assign N266 = in_sig[22] & \genblk2.roundPosMask [22];
  assign N268 = in_sig[21] & \genblk2.roundPosMask [21];
  assign N270 = in_sig[20] & \genblk2.roundPosMask [20];
  assign N272 = in_sig[19] & \genblk2.roundPosMask [19];
  assign N274 = in_sig[18] & \genblk2.roundPosMask [18];
  assign N276 = in_sig[17] & \genblk2.roundPosMask [17];
  assign N278 = in_sig[16] & \genblk2.roundPosMask [16];
  assign N280 = in_sig[15] & \genblk2.roundPosMask [15];
  assign N282 = in_sig[14] & \genblk2.roundPosMask [14];
  assign N284 = in_sig[13] & \genblk2.roundPosMask [13];
  assign N286 = in_sig[12] & \genblk2.roundPosMask [12];
  assign N288 = in_sig[11] & \genblk2.roundPosMask [11];
  assign N290 = in_sig[10] & \genblk2.roundPosMask [10];
  assign N292 = in_sig[9] & \genblk2.roundPosMask [9];
  assign N294 = in_sig[8] & \genblk2.roundPosMask [8];
  assign N296 = in_sig[7] & \genblk2.roundPosMask [7];
  assign N298 = in_sig[6] & \genblk2.roundPosMask [6];
  assign N300 = in_sig[5] & \genblk2.roundPosMask [5];
  assign N302 = in_sig[4] & \genblk2.roundPosMask [4];
  assign N304 = in_sig[3] & \genblk2.roundPosMask [3];
  assign N311 = N310 & N232;
  assign N310 = N308 | N309;
  assign N308 = N306 | N307;
  assign N306 = in_sig[2] & \genblk2.roundPosMask [2];
  assign N307 = in_sig[1] & \genblk2.roundPosMask [1];
  assign N309 = in_sig[0] & \genblk2.roundPosMask [0];
  assign \genblk2.anyRoundExtra  = N358 | N364;
  assign N358 = N356 | N357;
  assign N356 = N354 | N355;
  assign N354 = N352 | N353;
  assign N352 = N350 | N351;
  assign N350 = N348 | N349;
  assign N348 = N346 | N347;
  assign N346 = N344 | N345;
  assign N344 = N342 | N343;
  assign N342 = N340 | N341;
  assign N340 = N338 | N339;
  assign N338 = N336 | N337;
  assign N336 = N334 | N335;
  assign N334 = N332 | N333;
  assign N332 = N330 | N331;
  assign N330 = N328 | N329;
  assign N328 = N326 | N327;
  assign N326 = N324 | N325;
  assign N324 = N322 | N323;
  assign N322 = N320 | N321;
  assign N320 = N318 | N319;
  assign N318 = N316 | N317;
  assign N316 = N314 | N315;
  assign N314 = N312 | N313;
  assign N312 = in_sig[26] & 1'b0;
  assign N313 = in_sig[25] & \genblk2.genblk1.roundMask_main [24];
  assign N315 = in_sig[24] & \genblk2.genblk1.roundMask_main [23];
  assign N317 = in_sig[23] & \genblk2.genblk1.roundMask_main [22];
  assign N319 = in_sig[22] & \genblk2.genblk1.roundMask_main [21];
  assign N321 = in_sig[21] & \genblk2.genblk1.roundMask_main [20];
  assign N323 = in_sig[20] & \genblk2.genblk1.roundMask_main [19];
  assign N325 = in_sig[19] & \genblk2.genblk1.roundMask_main [18];
  assign N327 = in_sig[18] & \genblk2.genblk1.roundMask_main [17];
  assign N329 = in_sig[17] & \genblk2.genblk1.roundMask_main [16];
  assign N331 = in_sig[16] & \genblk2.genblk1.roundMask_main [15];
  assign N333 = in_sig[15] & \genblk2.genblk1.roundMask_main [14];
  assign N335 = in_sig[14] & \genblk2.genblk1.roundMask_main [13];
  assign N337 = in_sig[13] & \genblk2.genblk1.roundMask_main [12];
  assign N339 = in_sig[12] & \genblk2.genblk1.roundMask_main [11];
  assign N341 = in_sig[11] & \genblk2.genblk1.roundMask_main [10];
  assign N343 = in_sig[10] & \genblk2.genblk1.roundMask_main [9];
  assign N345 = in_sig[9] & \genblk2.genblk1.roundMask_main [8];
  assign N347 = in_sig[8] & \genblk2.genblk1.roundMask_main [7];
  assign N349 = in_sig[7] & \genblk2.genblk1.roundMask_main [6];
  assign N351 = in_sig[6] & \genblk2.genblk1.roundMask_main [5];
  assign N353 = in_sig[5] & \genblk2.genblk1.roundMask_main [4];
  assign N355 = in_sig[4] & \genblk2.genblk1.roundMask_main [3];
  assign N357 = in_sig[3] & \genblk2.genblk1.roundMask_main [2];
  assign N364 = N363 & N232;
  assign N363 = N361 | N362;
  assign N361 = N359 | N360;
  assign N359 = in_sig[2] & \genblk2.genblk1.roundMask_main [1];
  assign N360 = in_sig[1] & \genblk2.roundMask [2];
  assign N362 = in_sig[0] & 1'b1;
  assign \genblk2.anyRound  = \genblk2.roundPosBit  | \genblk2.anyRoundExtra ;
  assign \genblk2.roundIncr  = N366 | N367;
  assign N366 = N365 & \genblk2.roundPosBit ;
  assign N365 = N220 | N217;
  assign N367 = roundMagUp & \genblk2.anyRound ;
  assign N14 = ~\genblk2.roundIncr ;
  assign N15 = N368 & N369;
  assign N368 = N220 & \genblk2.roundPosBit ;
  assign N369 = ~\genblk2.anyRoundExtra ;
  assign N16 = ~N15;
  assign N42 = in_sig[26] | \genblk2.genblk1.roundMask_main [24];
  assign N43 = in_sig[25] | \genblk2.genblk1.roundMask_main [23];
  assign N44 = in_sig[24] | \genblk2.genblk1.roundMask_main [22];
  assign N45 = in_sig[23] | \genblk2.genblk1.roundMask_main [21];
  assign N46 = in_sig[22] | \genblk2.genblk1.roundMask_main [20];
  assign N47 = in_sig[21] | \genblk2.genblk1.roundMask_main [19];
  assign N48 = in_sig[20] | \genblk2.genblk1.roundMask_main [18];
  assign N49 = in_sig[19] | \genblk2.genblk1.roundMask_main [17];
  assign N50 = in_sig[18] | \genblk2.genblk1.roundMask_main [16];
  assign N51 = in_sig[17] | \genblk2.genblk1.roundMask_main [15];
  assign N52 = in_sig[16] | \genblk2.genblk1.roundMask_main [14];
  assign N53 = in_sig[15] | \genblk2.genblk1.roundMask_main [13];
  assign N54 = in_sig[14] | \genblk2.genblk1.roundMask_main [12];
  assign N55 = in_sig[13] | \genblk2.genblk1.roundMask_main [11];
  assign N56 = in_sig[12] | \genblk2.genblk1.roundMask_main [10];
  assign N57 = in_sig[11] | \genblk2.genblk1.roundMask_main [9];
  assign N58 = in_sig[10] | \genblk2.genblk1.roundMask_main [8];
  assign N59 = in_sig[9] | \genblk2.genblk1.roundMask_main [7];
  assign N60 = in_sig[8] | \genblk2.genblk1.roundMask_main [6];
  assign N61 = in_sig[7] | \genblk2.genblk1.roundMask_main [5];
  assign N62 = in_sig[6] | \genblk2.genblk1.roundMask_main [4];
  assign N63 = in_sig[5] | \genblk2.genblk1.roundMask_main [3];
  assign N64 = in_sig[4] | \genblk2.genblk1.roundMask_main [2];
  assign N65 = in_sig[3] | \genblk2.genblk1.roundMask_main [1];
  assign N66 = in_sig[2] | \genblk2.roundMask [2];
  assign N93 = N92 & N370;
  assign N370 = ~N41;
  assign N94 = N91 & N371;
  assign N371 = ~N40;
  assign N95 = N90 & N372;
  assign N372 = ~N39;
  assign N96 = N89 & N373;
  assign N373 = ~N38;
  assign N97 = N88 & N374;
  assign N374 = ~N37;
  assign N98 = N87 & N375;
  assign N375 = ~N36;
  assign N99 = N86 & N376;
  assign N376 = ~N35;
  assign N100 = N85 & N377;
  assign N377 = ~N34;
  assign N101 = N84 & N378;
  assign N378 = ~N33;
  assign N102 = N83 & N379;
  assign N379 = ~N32;
  assign N103 = N82 & N380;
  assign N380 = ~N31;
  assign N104 = N81 & N381;
  assign N381 = ~N30;
  assign N105 = N80 & N382;
  assign N382 = ~N29;
  assign N106 = N79 & N383;
  assign N383 = ~N28;
  assign N107 = N78 & N384;
  assign N384 = ~N27;
  assign N108 = N77 & N385;
  assign N385 = ~N26;
  assign N109 = N76 & N386;
  assign N386 = ~N25;
  assign N110 = N75 & N387;
  assign N387 = ~N24;
  assign N111 = N74 & N388;
  assign N388 = ~N23;
  assign N112 = N73 & N389;
  assign N389 = ~N22;
  assign N113 = N72 & N390;
  assign N390 = ~N21;
  assign N114 = N71 & N391;
  assign N391 = ~N20;
  assign N115 = N70 & N392;
  assign N392 = ~N19;
  assign N116 = N69 & N393;
  assign N393 = ~N18;
  assign N117 = N68 & N394;
  assign N394 = ~N17;
  assign N118 = N67 & N395;
  assign N395 = ~N15;
  assign N119 = N214 & \genblk2.anyRound ;
  assign N120 = ~N119;
  assign N147 = N396 | N145;
  assign N396 = in_sig[26] & N233;
  assign N148 = N397 | N144;
  assign N397 = in_sig[25] & N234;
  assign N149 = N398 | N143;
  assign N398 = in_sig[24] & N235;
  assign N150 = N399 | N142;
  assign N399 = in_sig[23] & N236;
  assign N151 = N400 | N141;
  assign N400 = in_sig[22] & N237;
  assign N152 = N401 | N140;
  assign N401 = in_sig[21] & N238;
  assign N153 = N402 | N139;
  assign N402 = in_sig[20] & N239;
  assign N154 = N403 | N138;
  assign N403 = in_sig[19] & N240;
  assign N155 = N404 | N137;
  assign N404 = in_sig[18] & N241;
  assign N156 = N405 | N136;
  assign N405 = in_sig[17] & N242;
  assign N157 = N406 | N135;
  assign N406 = in_sig[16] & N243;
  assign N158 = N407 | N134;
  assign N407 = in_sig[15] & N244;
  assign N159 = N408 | N133;
  assign N408 = in_sig[14] & N245;
  assign N160 = N409 | N132;
  assign N409 = in_sig[13] & N246;
  assign N161 = N410 | N131;
  assign N410 = in_sig[12] & N247;
  assign N162 = N411 | N130;
  assign N411 = in_sig[11] & N248;
  assign N163 = N412 | N129;
  assign N412 = in_sig[10] & N249;
  assign N164 = N413 | N128;
  assign N413 = in_sig[9] & N250;
  assign N165 = N414 | N127;
  assign N414 = in_sig[8] & N251;
  assign N166 = N415 | N126;
  assign N415 = in_sig[7] & N252;
  assign N167 = N416 | N125;
  assign N416 = in_sig[6] & N253;
  assign N168 = N417 | N124;
  assign N417 = in_sig[5] & N254;
  assign N169 = N418 | N123;
  assign N418 = in_sig[4] & N255;
  assign N170 = N419 | N122;
  assign N419 = in_sig[3] & N256;
  assign N171 = N420 | N121;
  assign N420 = in_sig[2] & N257;
  assign N172 = ~in_sig[26];
  assign \genblk2.unboundedRange_anyRound  = N421 | N422;
  assign N421 = in_sig[26] & in_sig[2];
  assign N422 = in_sig[1] | in_sig[0];
  assign \genblk2.unboundedRange_roundIncr  = N424 | N425;
  assign N424 = N423 & \genblk2.unboundedRange_roundPosBit ;
  assign N423 = N220 | N217;
  assign N425 = roundMagUp & \genblk2.unboundedRange_anyRound ;
  assign N175 = \genblk2.anyRound  & N174;
  assign N176 = ~N175;
  assign N179 = ~control[0];
  assign N180 = ~N178;
  assign common_underflow = common_totalUnderflow | N430;
  assign N430 = N177 & N429;
  assign N429 = ~N428;
  assign N428 = N427 & \genblk2.unboundedRange_roundIncr ;
  assign N427 = N426 & \genblk2.roundPosBit ;
  assign N426 = N181 & \genblk2.roundCarry ;
  assign common_inexact = common_totalUnderflow | \genblk2.anyRound ;
  assign notNaN_isSpecialInfOut = exceptionFlags_3_ | in_isInf;
  assign commonCase = N433 & N434;
  assign N433 = N431 & N432;
  assign N431 = ~isNaNOut;
  assign N432 = ~notNaN_isSpecialInfOut;
  assign N434 = ~in_isZero;
  assign exceptionFlags[2] = commonCase & common_overflow;
  assign exceptionFlags[1] = commonCase & common_underflow;
  assign exceptionFlags[0] = exceptionFlags[2] | N435;
  assign N435 = commonCase & common_inexact;
  assign overflow_roundMagUp = N436 | roundMagUp;
  assign N436 = N220 | N217;
  assign pegMinNonzeroMagOut = N437 & N438;
  assign N437 = commonCase & common_totalUnderflow;
  assign N438 = roundMagUp | N214;
  assign pegMaxFiniteMagOut = exceptionFlags[2] & N439;
  assign N439 = ~overflow_roundMagUp;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | N440;
  assign N440 = exceptionFlags[2] & overflow_roundMagUp;
  assign N182 = in_isZero | common_totalUnderflow;
  assign out[31] = N446 | isNaNOut;
  assign N446 = N445 | notNaN_isInfOut;
  assign N445 = N444 | pegMaxFiniteMagOut;
  assign N444 = N442 & N443;
  assign N442 = \genblk2.sRoundedExp [8] & N441;
  assign N441 = ~N182;
  assign N443 = ~pegMinNonzeroMagOut;
  assign out[30] = N451 | isNaNOut;
  assign N451 = N450 | notNaN_isInfOut;
  assign N450 = N448 & N449;
  assign N448 = N447 & N443;
  assign N447 = \genblk2.sRoundedExp [7] & N441;
  assign N449 = ~pegMaxFiniteMagOut;
  assign out[29] = N456 | isNaNOut;
  assign N456 = N455 | pegMaxFiniteMagOut;
  assign N455 = N454 | pegMinNonzeroMagOut;
  assign N454 = N452 & N453;
  assign N452 = \genblk2.sRoundedExp [6] & N441;
  assign N453 = ~notNaN_isInfOut;
  assign out[28] = N457 | pegMaxFiniteMagOut;
  assign N457 = \genblk2.sRoundedExp [5] | pegMinNonzeroMagOut;
  assign out[27] = N458 | pegMaxFiniteMagOut;
  assign N458 = \genblk2.sRoundedExp [4] & N443;
  assign out[26] = N459 | pegMaxFiniteMagOut;
  assign N459 = \genblk2.sRoundedExp [3] | pegMinNonzeroMagOut;
  assign out[25] = N460 | pegMaxFiniteMagOut;
  assign N460 = \genblk2.sRoundedExp [2] & N443;
  assign out[24] = N461 | pegMaxFiniteMagOut;
  assign N461 = \genblk2.sRoundedExp [1] | pegMinNonzeroMagOut;
  assign out[23] = N462 | pegMaxFiniteMagOut;
  assign N462 = \genblk2.sRoundedExp [0] | pegMinNonzeroMagOut;
  assign N183 = N434 & N463;
  assign N463 = ~common_totalUnderflow;
  assign N184 = ~N183;
  assign N186 = N464 & N463;
  assign N464 = N431 & N434;
  assign N187 = ~N186;
  assign out[22] = N465 | pegMaxFiniteMagOut;
  assign N465 = isNaNOut | N185;
  assign out[21] = N209 | pegMaxFiniteMagOut;
  assign out[20] = N208 | pegMaxFiniteMagOut;
  assign out[19] = N207 | pegMaxFiniteMagOut;
  assign out[18] = N206 | pegMaxFiniteMagOut;
  assign out[17] = N205 | pegMaxFiniteMagOut;
  assign out[16] = N204 | pegMaxFiniteMagOut;
  assign out[15] = N203 | pegMaxFiniteMagOut;
  assign out[14] = N202 | pegMaxFiniteMagOut;
  assign out[13] = N201 | pegMaxFiniteMagOut;
  assign out[12] = N200 | pegMaxFiniteMagOut;
  assign out[11] = N199 | pegMaxFiniteMagOut;
  assign out[10] = N198 | pegMaxFiniteMagOut;
  assign out[9] = N197 | pegMaxFiniteMagOut;
  assign out[8] = N196 | pegMaxFiniteMagOut;
  assign out[7] = N195 | pegMaxFiniteMagOut;
  assign out[6] = N194 | pegMaxFiniteMagOut;
  assign out[5] = N193 | pegMaxFiniteMagOut;
  assign out[4] = N192 | pegMaxFiniteMagOut;
  assign out[3] = N191 | pegMaxFiniteMagOut;
  assign out[2] = N190 | pegMaxFiniteMagOut;
  assign out[1] = N189 | pegMaxFiniteMagOut;
  assign out[0] = N188 | pegMaxFiniteMagOut;

endmodule



module roundRawFNToRecFN_expWidth8_sigWidth24
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [9:0] in_sExp;
  input [26:0] in_sig;
  input [2:0] roundingMode;
  output [32:0] out;
  output [4:0] exceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [32:0] out;
  wire [4:0] exceptionFlags;

  roundAnyRawFNToRecFN_inExpWidth8_inSigWidth26_outExpWidth8_outSigWidth24_options0
  roundAnyRawFNToRecFN
  (
    .control(control[0]),
    .invalidExc(invalidExc),
    .infiniteExc(infiniteExc),
    .in_isNaN(in_isNaN),
    .in_isInf(in_isInf),
    .in_isZero(in_isZero),
    .in_sign(in_sign),
    .in_sExp(in_sExp),
    .in_sig(in_sig),
    .roundingMode(roundingMode),
    .out(out),
    .exceptionFlags(exceptionFlags)
  );


endmodule



module fpu_float_fma_round
(
  clk_i,
  reset_i,
  stall_fpu2_i,
  fma1_v_i,
  fma1_rm_i,
  invalidExc_i,
  in_isNaN_i,
  in_isInf_i,
  in_isZero_i,
  in_sign_i,
  in_sExp_i,
  in_sig_i,
  fma2_v_o,
  fma2_result_o,
  fma2_fflags_o_invalid_,
  fma2_fflags_o_div_zero_,
  fma2_fflags_o_overflow_,
  fma2_fflags_o_underflow_,
  fma2_fflags_o_inexact_
);

  input [2:0] fma1_rm_i;
  input [9:0] in_sExp_i;
  input [26:0] in_sig_i;
  output [32:0] fma2_result_o;
  input clk_i;
  input reset_i;
  input stall_fpu2_i;
  input fma1_v_i;
  input invalidExc_i;
  input in_isNaN_i;
  input in_isInf_i;
  input in_isZero_i;
  input in_sign_i;
  output fma2_v_o;
  output fma2_fflags_o_invalid_;
  output fma2_fflags_o_div_zero_;
  output fma2_fflags_o_overflow_;
  output fma2_fflags_o_underflow_;
  output fma2_fflags_o_inexact_;
  wire [32:0] fma2_result_o,result_lo;
  wire fma2_v_o,fma2_fflags_o_invalid_,fma2_fflags_o_div_zero_,fma2_fflags_o_overflow_,
  fma2_fflags_o_underflow_,fma2_fflags_o_inexact_,N0,N1,N3,fflags_lo_invalid_,
  fflags_lo_div_zero_,fflags_lo_overflow_,fflags_lo_underflow_,fflags_lo_inexact_,N4,
  N5,N6,N7,N8,N9,N10;
  reg fma2_result_o_32_sv2v_reg,fma2_result_o_31_sv2v_reg,fma2_result_o_30_sv2v_reg,
  fma2_result_o_29_sv2v_reg,fma2_result_o_28_sv2v_reg,fma2_result_o_27_sv2v_reg,
  fma2_result_o_26_sv2v_reg,fma2_result_o_25_sv2v_reg,fma2_result_o_24_sv2v_reg,
  fma2_result_o_23_sv2v_reg,fma2_result_o_22_sv2v_reg,fma2_result_o_21_sv2v_reg,
  fma2_result_o_20_sv2v_reg,fma2_result_o_19_sv2v_reg,fma2_result_o_18_sv2v_reg,
  fma2_result_o_17_sv2v_reg,fma2_result_o_16_sv2v_reg,fma2_result_o_15_sv2v_reg,
  fma2_result_o_14_sv2v_reg,fma2_result_o_13_sv2v_reg,fma2_result_o_12_sv2v_reg,
  fma2_result_o_11_sv2v_reg,fma2_result_o_10_sv2v_reg,fma2_result_o_9_sv2v_reg,
  fma2_result_o_8_sv2v_reg,fma2_result_o_7_sv2v_reg,fma2_result_o_6_sv2v_reg,
  fma2_result_o_5_sv2v_reg,fma2_result_o_4_sv2v_reg,fma2_result_o_3_sv2v_reg,fma2_result_o_2_sv2v_reg,
  fma2_result_o_1_sv2v_reg,fma2_result_o_0_sv2v_reg,fma2_v_o_sv2v_reg,
  fma2_fflags_o_invalid__sv2v_reg,fma2_fflags_o_div_zero__sv2v_reg,
  fma2_fflags_o_overflow__sv2v_reg,fma2_fflags_o_underflow__sv2v_reg,fma2_fflags_o_inexact__sv2v_reg;
  assign fma2_result_o[32] = fma2_result_o_32_sv2v_reg;
  assign fma2_result_o[31] = fma2_result_o_31_sv2v_reg;
  assign fma2_result_o[30] = fma2_result_o_30_sv2v_reg;
  assign fma2_result_o[29] = fma2_result_o_29_sv2v_reg;
  assign fma2_result_o[28] = fma2_result_o_28_sv2v_reg;
  assign fma2_result_o[27] = fma2_result_o_27_sv2v_reg;
  assign fma2_result_o[26] = fma2_result_o_26_sv2v_reg;
  assign fma2_result_o[25] = fma2_result_o_25_sv2v_reg;
  assign fma2_result_o[24] = fma2_result_o_24_sv2v_reg;
  assign fma2_result_o[23] = fma2_result_o_23_sv2v_reg;
  assign fma2_result_o[22] = fma2_result_o_22_sv2v_reg;
  assign fma2_result_o[21] = fma2_result_o_21_sv2v_reg;
  assign fma2_result_o[20] = fma2_result_o_20_sv2v_reg;
  assign fma2_result_o[19] = fma2_result_o_19_sv2v_reg;
  assign fma2_result_o[18] = fma2_result_o_18_sv2v_reg;
  assign fma2_result_o[17] = fma2_result_o_17_sv2v_reg;
  assign fma2_result_o[16] = fma2_result_o_16_sv2v_reg;
  assign fma2_result_o[15] = fma2_result_o_15_sv2v_reg;
  assign fma2_result_o[14] = fma2_result_o_14_sv2v_reg;
  assign fma2_result_o[13] = fma2_result_o_13_sv2v_reg;
  assign fma2_result_o[12] = fma2_result_o_12_sv2v_reg;
  assign fma2_result_o[11] = fma2_result_o_11_sv2v_reg;
  assign fma2_result_o[10] = fma2_result_o_10_sv2v_reg;
  assign fma2_result_o[9] = fma2_result_o_9_sv2v_reg;
  assign fma2_result_o[8] = fma2_result_o_8_sv2v_reg;
  assign fma2_result_o[7] = fma2_result_o_7_sv2v_reg;
  assign fma2_result_o[6] = fma2_result_o_6_sv2v_reg;
  assign fma2_result_o[5] = fma2_result_o_5_sv2v_reg;
  assign fma2_result_o[4] = fma2_result_o_4_sv2v_reg;
  assign fma2_result_o[3] = fma2_result_o_3_sv2v_reg;
  assign fma2_result_o[2] = fma2_result_o_2_sv2v_reg;
  assign fma2_result_o[1] = fma2_result_o_1_sv2v_reg;
  assign fma2_result_o[0] = fma2_result_o_0_sv2v_reg;
  assign fma2_v_o = fma2_v_o_sv2v_reg;
  assign fma2_fflags_o_invalid_ = fma2_fflags_o_invalid__sv2v_reg;
  assign fma2_fflags_o_div_zero_ = fma2_fflags_o_div_zero__sv2v_reg;
  assign fma2_fflags_o_overflow_ = fma2_fflags_o_overflow__sv2v_reg;
  assign fma2_fflags_o_underflow_ = fma2_fflags_o_underflow__sv2v_reg;
  assign fma2_fflags_o_inexact_ = fma2_fflags_o_inexact__sv2v_reg;

  roundRawFNToRecFN_expWidth8_sigWidth24
  round0
  (
    .control(1'b1),
    .invalidExc(invalidExc_i),
    .infiniteExc(1'b0),
    .in_isNaN(in_isNaN_i),
    .in_isInf(in_isInf_i),
    .in_isZero(in_isZero_i),
    .in_sign(in_sign_i),
    .in_sExp(in_sExp_i),
    .in_sig(in_sig_i),
    .roundingMode(fma1_rm_i),
    .out(result_lo),
    .exceptionFlags({ fflags_lo_invalid_, fflags_lo_div_zero_, fflags_lo_overflow_, fflags_lo_underflow_, fflags_lo_inexact_ })
  );

  assign N7 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = N4;
  assign N1 = stall_fpu2_i;
  assign N8 = (N3)? 1'b0 : 
              (N10)? fma1_v_i : 
              (N6)? 1'b0 : 1'b0;
  assign N3 = reset_i;
  assign N4 = ~stall_fpu2_i;
  assign N5 = N4 | reset_i;
  assign N6 = ~N5;
  assign N9 = ~reset_i;
  assign N10 = N4 & N9;

  always @(posedge clk_i) begin
    if(N8) begin
      fma2_result_o_32_sv2v_reg <= result_lo[32];
      fma2_result_o_31_sv2v_reg <= result_lo[31];
      fma2_result_o_30_sv2v_reg <= result_lo[30];
      fma2_result_o_29_sv2v_reg <= result_lo[29];
      fma2_result_o_28_sv2v_reg <= result_lo[28];
      fma2_result_o_27_sv2v_reg <= result_lo[27];
      fma2_result_o_26_sv2v_reg <= result_lo[26];
      fma2_result_o_25_sv2v_reg <= result_lo[25];
      fma2_result_o_24_sv2v_reg <= result_lo[24];
      fma2_result_o_23_sv2v_reg <= result_lo[23];
      fma2_result_o_22_sv2v_reg <= result_lo[22];
      fma2_result_o_21_sv2v_reg <= result_lo[21];
      fma2_result_o_20_sv2v_reg <= result_lo[20];
      fma2_result_o_19_sv2v_reg <= result_lo[19];
      fma2_result_o_18_sv2v_reg <= result_lo[18];
      fma2_result_o_17_sv2v_reg <= result_lo[17];
      fma2_result_o_16_sv2v_reg <= result_lo[16];
      fma2_result_o_15_sv2v_reg <= result_lo[15];
      fma2_result_o_14_sv2v_reg <= result_lo[14];
      fma2_result_o_13_sv2v_reg <= result_lo[13];
      fma2_result_o_12_sv2v_reg <= result_lo[12];
      fma2_result_o_11_sv2v_reg <= result_lo[11];
      fma2_result_o_10_sv2v_reg <= result_lo[10];
      fma2_result_o_9_sv2v_reg <= result_lo[9];
      fma2_result_o_8_sv2v_reg <= result_lo[8];
      fma2_result_o_7_sv2v_reg <= result_lo[7];
      fma2_result_o_6_sv2v_reg <= result_lo[6];
      fma2_result_o_5_sv2v_reg <= result_lo[5];
      fma2_result_o_4_sv2v_reg <= result_lo[4];
      fma2_result_o_3_sv2v_reg <= result_lo[3];
      fma2_result_o_2_sv2v_reg <= result_lo[2];
      fma2_result_o_1_sv2v_reg <= result_lo[1];
      fma2_result_o_0_sv2v_reg <= result_lo[0];
      fma2_fflags_o_invalid__sv2v_reg <= fflags_lo_invalid_;
      fma2_fflags_o_div_zero__sv2v_reg <= fflags_lo_div_zero_;
      fma2_fflags_o_overflow__sv2v_reg <= fflags_lo_overflow_;
      fma2_fflags_o_underflow__sv2v_reg <= fflags_lo_underflow_;
      fma2_fflags_o_inexact__sv2v_reg <= fflags_lo_inexact_;
    end 
    if(reset_i) begin
      fma2_v_o_sv2v_reg <= 1'b0;
    end else if(N7) begin
      fma2_v_o_sv2v_reg <= fma1_v_i;
    end 
  end


endmodule



module reverse_width32
(
  in,
  out
);

  input [31:0] in;
  output [31:0] out;
  wire [31:0] out;
  assign out[31] = in[0];
  assign out[30] = in[1];
  assign out[29] = in[2];
  assign out[28] = in[3];
  assign out[27] = in[4];
  assign out[26] = in[5];
  assign out[25] = in[6];
  assign out[24] = in[7];
  assign out[23] = in[8];
  assign out[22] = in[9];
  assign out[21] = in[10];
  assign out[20] = in[11];
  assign out[19] = in[12];
  assign out[18] = in[13];
  assign out[17] = in[14];
  assign out[16] = in[15];
  assign out[15] = in[16];
  assign out[14] = in[17];
  assign out[13] = in[18];
  assign out[12] = in[19];
  assign out[11] = in[20];
  assign out[10] = in[21];
  assign out[9] = in[22];
  assign out[8] = in[23];
  assign out[7] = in[24];
  assign out[6] = in[25];
  assign out[5] = in[26];
  assign out[4] = in[27];
  assign out[3] = in[28];
  assign out[2] = in[29];
  assign out[1] = in[30];
  assign out[0] = in[31];

endmodule



module countLeadingZeros_inWidth32_countWidth5
(
  in,
  count
);

  input [31:0] in;
  output [4:0] count;
  wire [4:0] count;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,\Bit_5_.countSoFar_0 ,\Bit_9_.countSoFar_0 ,\Bit_10_.countSoFar_1 ,
  \Bit_11_.countSoFar_3 ,\Bit_13_.countSoFar_0 ,\Bit_17_.countSoFar_0 ,
  \Bit_18_.countSoFar_1 ,\Bit_19_.countSoFar_4 ,\Bit_20_.countSoFar_2 ,\Bit_21_.countSoFar_2 ,
  \Bit_21_.countSoFar_0 ,\Bit_22_.countSoFar_4 ,\Bit_23_.countSoFar_4 ,
  \Bit_25_.countSoFar_0 ,\Bit_26_.countSoFar_1 ,\Bit_27_.countSoFar_1 ,\Bit_27_.countSoFar_0 ,
  \Bit_29_.countSoFar_0 ,sv2v_dc_1;
  wire [31:0] reverseIn;
  wire [31:1] oneLeastReverseIn;
  wire [0:0] \Bit_1_.countSoFar ;
  wire [1:1] \Bit_2_.countSoFar ;
  wire [1:0] \Bit_3_.countSoFar ,\Bit_11_.countSoFar ,\Bit_19_.countSoFar ;
  wire [2:2] \Bit_4_.countSoFar ,\Bit_5_.countSoFar ;
  wire [2:1] \Bit_6_.countSoFar ,\Bit_22_.countSoFar ;
  wire [2:0] \Bit_7_.countSoFar ,\Bit_23_.countSoFar ;
  wire [3:3] \Bit_8_.countSoFar ,\Bit_9_.countSoFar ,\Bit_10_.countSoFar ;
  wire [3:2] \Bit_12_.countSoFar ,\Bit_13_.countSoFar ;
  wire [3:1] \Bit_14_.countSoFar ;
  wire [3:0] \Bit_15_.countSoFar ;
  wire [4:4] \Bit_16_.countSoFar ,\Bit_17_.countSoFar ,\Bit_18_.countSoFar ,
  \Bit_20_.countSoFar ,\Bit_21_.countSoFar ;
  wire [4:3] \Bit_24_.countSoFar ,\Bit_25_.countSoFar ,\Bit_26_.countSoFar ,
  \Bit_27_.countSoFar ;
  wire [4:2] \Bit_28_.countSoFar ,\Bit_29_.countSoFar ;
  wire [4:1] \Bit_30_.countSoFar ;

  reverse_width32
  reverse_in
  (
    .in(in),
    .out(reverseIn)
  );

  assign { N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, sv2v_dc_1 } = { N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31 } + 1'b1;
  assign N0 = ~reverseIn[31];
  assign N1 = ~reverseIn[30];
  assign N2 = ~reverseIn[29];
  assign N3 = ~reverseIn[28];
  assign N4 = ~reverseIn[27];
  assign N5 = ~reverseIn[26];
  assign N6 = ~reverseIn[25];
  assign N7 = ~reverseIn[24];
  assign N8 = ~reverseIn[23];
  assign N9 = ~reverseIn[22];
  assign N10 = ~reverseIn[21];
  assign N11 = ~reverseIn[20];
  assign N12 = ~reverseIn[19];
  assign N13 = ~reverseIn[18];
  assign N14 = ~reverseIn[17];
  assign N15 = ~reverseIn[16];
  assign N16 = ~reverseIn[15];
  assign N17 = ~reverseIn[14];
  assign N18 = ~reverseIn[13];
  assign N19 = ~reverseIn[12];
  assign N20 = ~reverseIn[11];
  assign N21 = ~reverseIn[10];
  assign N22 = ~reverseIn[9];
  assign N23 = ~reverseIn[8];
  assign N24 = ~reverseIn[7];
  assign N25 = ~reverseIn[6];
  assign N26 = ~reverseIn[5];
  assign N27 = ~reverseIn[4];
  assign N28 = ~reverseIn[3];
  assign N29 = ~reverseIn[2];
  assign N30 = ~reverseIn[1];
  assign N31 = ~reverseIn[0];
  assign oneLeastReverseIn[31] = reverseIn[31] & N62;
  assign oneLeastReverseIn[30] = reverseIn[30] & N61;
  assign oneLeastReverseIn[29] = reverseIn[29] & N60;
  assign oneLeastReverseIn[28] = reverseIn[28] & N59;
  assign oneLeastReverseIn[27] = reverseIn[27] & N58;
  assign oneLeastReverseIn[26] = reverseIn[26] & N57;
  assign oneLeastReverseIn[25] = reverseIn[25] & N56;
  assign oneLeastReverseIn[24] = reverseIn[24] & N55;
  assign oneLeastReverseIn[23] = reverseIn[23] & N54;
  assign oneLeastReverseIn[22] = reverseIn[22] & N53;
  assign oneLeastReverseIn[21] = reverseIn[21] & N52;
  assign oneLeastReverseIn[20] = reverseIn[20] & N51;
  assign oneLeastReverseIn[19] = reverseIn[19] & N50;
  assign oneLeastReverseIn[18] = reverseIn[18] & N49;
  assign oneLeastReverseIn[17] = reverseIn[17] & N48;
  assign oneLeastReverseIn[16] = reverseIn[16] & N47;
  assign oneLeastReverseIn[15] = reverseIn[15] & N46;
  assign oneLeastReverseIn[14] = reverseIn[14] & N45;
  assign oneLeastReverseIn[13] = reverseIn[13] & N44;
  assign oneLeastReverseIn[12] = reverseIn[12] & N43;
  assign oneLeastReverseIn[11] = reverseIn[11] & N42;
  assign oneLeastReverseIn[10] = reverseIn[10] & N41;
  assign oneLeastReverseIn[9] = reverseIn[9] & N40;
  assign oneLeastReverseIn[8] = reverseIn[8] & N39;
  assign oneLeastReverseIn[7] = reverseIn[7] & N38;
  assign oneLeastReverseIn[6] = reverseIn[6] & N37;
  assign oneLeastReverseIn[5] = reverseIn[5] & N36;
  assign oneLeastReverseIn[4] = reverseIn[4] & N35;
  assign oneLeastReverseIn[3] = reverseIn[3] & N34;
  assign oneLeastReverseIn[2] = reverseIn[2] & N33;
  assign oneLeastReverseIn[1] = reverseIn[1] & N32;
  assign \Bit_1_.countSoFar [0] = 1'b0 | oneLeastReverseIn[1];
  assign \Bit_2_.countSoFar [1] = 1'b0 | oneLeastReverseIn[2];
  assign \Bit_3_.countSoFar [1] = \Bit_2_.countSoFar [1] | oneLeastReverseIn[3];
  assign \Bit_3_.countSoFar [0] = \Bit_1_.countSoFar [0] | oneLeastReverseIn[3];
  assign \Bit_4_.countSoFar [2] = 1'b0 | oneLeastReverseIn[4];
  assign \Bit_5_.countSoFar [2] = \Bit_4_.countSoFar [2] | oneLeastReverseIn[5];
  assign \Bit_5_.countSoFar_0  = \Bit_3_.countSoFar [0] | oneLeastReverseIn[5];
  assign \Bit_6_.countSoFar [2] = \Bit_5_.countSoFar [2] | oneLeastReverseIn[6];
  assign \Bit_6_.countSoFar [1] = \Bit_3_.countSoFar [1] | oneLeastReverseIn[6];
  assign \Bit_7_.countSoFar [2] = \Bit_6_.countSoFar [2] | oneLeastReverseIn[7];
  assign \Bit_7_.countSoFar [1] = \Bit_6_.countSoFar [1] | oneLeastReverseIn[7];
  assign \Bit_7_.countSoFar [0] = \Bit_5_.countSoFar_0  | oneLeastReverseIn[7];
  assign \Bit_8_.countSoFar [3] = 1'b0 | oneLeastReverseIn[8];
  assign \Bit_9_.countSoFar [3] = \Bit_8_.countSoFar [3] | oneLeastReverseIn[9];
  assign \Bit_9_.countSoFar_0  = \Bit_7_.countSoFar [0] | oneLeastReverseIn[9];
  assign \Bit_10_.countSoFar [3] = \Bit_9_.countSoFar [3] | oneLeastReverseIn[10];
  assign \Bit_10_.countSoFar_1  = \Bit_7_.countSoFar [1] | oneLeastReverseIn[10];
  assign \Bit_11_.countSoFar_3  = \Bit_10_.countSoFar [3] | oneLeastReverseIn[11];
  assign \Bit_11_.countSoFar [1] = \Bit_10_.countSoFar_1  | oneLeastReverseIn[11];
  assign \Bit_11_.countSoFar [0] = \Bit_9_.countSoFar_0  | oneLeastReverseIn[11];
  assign \Bit_12_.countSoFar [3] = \Bit_11_.countSoFar_3  | oneLeastReverseIn[12];
  assign \Bit_12_.countSoFar [2] = \Bit_7_.countSoFar [2] | oneLeastReverseIn[12];
  assign \Bit_13_.countSoFar [3] = \Bit_12_.countSoFar [3] | oneLeastReverseIn[13];
  assign \Bit_13_.countSoFar [2] = \Bit_12_.countSoFar [2] | oneLeastReverseIn[13];
  assign \Bit_13_.countSoFar_0  = \Bit_11_.countSoFar [0] | oneLeastReverseIn[13];
  assign \Bit_14_.countSoFar [3] = \Bit_13_.countSoFar [3] | oneLeastReverseIn[14];
  assign \Bit_14_.countSoFar [2] = \Bit_13_.countSoFar [2] | oneLeastReverseIn[14];
  assign \Bit_14_.countSoFar [1] = \Bit_11_.countSoFar [1] | oneLeastReverseIn[14];
  assign \Bit_15_.countSoFar [3] = \Bit_14_.countSoFar [3] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [2] = \Bit_14_.countSoFar [2] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [1] = \Bit_14_.countSoFar [1] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [0] = \Bit_13_.countSoFar_0  | oneLeastReverseIn[15];
  assign \Bit_16_.countSoFar [4] = 1'b0 | oneLeastReverseIn[16];
  assign \Bit_17_.countSoFar [4] = \Bit_16_.countSoFar [4] | oneLeastReverseIn[17];
  assign \Bit_17_.countSoFar_0  = \Bit_15_.countSoFar [0] | oneLeastReverseIn[17];
  assign \Bit_18_.countSoFar [4] = \Bit_17_.countSoFar [4] | oneLeastReverseIn[18];
  assign \Bit_18_.countSoFar_1  = \Bit_15_.countSoFar [1] | oneLeastReverseIn[18];
  assign \Bit_19_.countSoFar_4  = \Bit_18_.countSoFar [4] | oneLeastReverseIn[19];
  assign \Bit_19_.countSoFar [1] = \Bit_18_.countSoFar_1  | oneLeastReverseIn[19];
  assign \Bit_19_.countSoFar [0] = \Bit_17_.countSoFar_0  | oneLeastReverseIn[19];
  assign \Bit_20_.countSoFar [4] = \Bit_19_.countSoFar_4  | oneLeastReverseIn[20];
  assign \Bit_20_.countSoFar_2  = \Bit_15_.countSoFar [2] | oneLeastReverseIn[20];
  assign \Bit_21_.countSoFar [4] = \Bit_20_.countSoFar [4] | oneLeastReverseIn[21];
  assign \Bit_21_.countSoFar_2  = \Bit_20_.countSoFar_2  | oneLeastReverseIn[21];
  assign \Bit_21_.countSoFar_0  = \Bit_19_.countSoFar [0] | oneLeastReverseIn[21];
  assign \Bit_22_.countSoFar_4  = \Bit_21_.countSoFar [4] | oneLeastReverseIn[22];
  assign \Bit_22_.countSoFar [2] = \Bit_21_.countSoFar_2  | oneLeastReverseIn[22];
  assign \Bit_22_.countSoFar [1] = \Bit_19_.countSoFar [1] | oneLeastReverseIn[22];
  assign \Bit_23_.countSoFar_4  = \Bit_22_.countSoFar_4  | oneLeastReverseIn[23];
  assign \Bit_23_.countSoFar [2] = \Bit_22_.countSoFar [2] | oneLeastReverseIn[23];
  assign \Bit_23_.countSoFar [1] = \Bit_22_.countSoFar [1] | oneLeastReverseIn[23];
  assign \Bit_23_.countSoFar [0] = \Bit_21_.countSoFar_0  | oneLeastReverseIn[23];
  assign \Bit_24_.countSoFar [4] = \Bit_23_.countSoFar_4  | oneLeastReverseIn[24];
  assign \Bit_24_.countSoFar [3] = \Bit_15_.countSoFar [3] | oneLeastReverseIn[24];
  assign \Bit_25_.countSoFar [4] = \Bit_24_.countSoFar [4] | oneLeastReverseIn[25];
  assign \Bit_25_.countSoFar [3] = \Bit_24_.countSoFar [3] | oneLeastReverseIn[25];
  assign \Bit_25_.countSoFar_0  = \Bit_23_.countSoFar [0] | oneLeastReverseIn[25];
  assign \Bit_26_.countSoFar [4] = \Bit_25_.countSoFar [4] | oneLeastReverseIn[26];
  assign \Bit_26_.countSoFar [3] = \Bit_25_.countSoFar [3] | oneLeastReverseIn[26];
  assign \Bit_26_.countSoFar_1  = \Bit_23_.countSoFar [1] | oneLeastReverseIn[26];
  assign \Bit_27_.countSoFar [4] = \Bit_26_.countSoFar [4] | oneLeastReverseIn[27];
  assign \Bit_27_.countSoFar [3] = \Bit_26_.countSoFar [3] | oneLeastReverseIn[27];
  assign \Bit_27_.countSoFar_1  = \Bit_26_.countSoFar_1  | oneLeastReverseIn[27];
  assign \Bit_27_.countSoFar_0  = \Bit_25_.countSoFar_0  | oneLeastReverseIn[27];
  assign \Bit_28_.countSoFar [4] = \Bit_27_.countSoFar [4] | oneLeastReverseIn[28];
  assign \Bit_28_.countSoFar [3] = \Bit_27_.countSoFar [3] | oneLeastReverseIn[28];
  assign \Bit_28_.countSoFar [2] = \Bit_23_.countSoFar [2] | oneLeastReverseIn[28];
  assign \Bit_29_.countSoFar [4] = \Bit_28_.countSoFar [4] | oneLeastReverseIn[29];
  assign \Bit_29_.countSoFar [3] = \Bit_28_.countSoFar [3] | oneLeastReverseIn[29];
  assign \Bit_29_.countSoFar [2] = \Bit_28_.countSoFar [2] | oneLeastReverseIn[29];
  assign \Bit_29_.countSoFar_0  = \Bit_27_.countSoFar_0  | oneLeastReverseIn[29];
  assign \Bit_30_.countSoFar [4] = \Bit_29_.countSoFar [4] | oneLeastReverseIn[30];
  assign \Bit_30_.countSoFar [3] = \Bit_29_.countSoFar [3] | oneLeastReverseIn[30];
  assign \Bit_30_.countSoFar [2] = \Bit_29_.countSoFar [2] | oneLeastReverseIn[30];
  assign \Bit_30_.countSoFar [1] = \Bit_27_.countSoFar_1  | oneLeastReverseIn[30];
  assign count[4] = \Bit_30_.countSoFar [4] | oneLeastReverseIn[31];
  assign count[3] = \Bit_30_.countSoFar [3] | oneLeastReverseIn[31];
  assign count[2] = \Bit_30_.countSoFar [2] | oneLeastReverseIn[31];
  assign count[1] = \Bit_30_.countSoFar [1] | oneLeastReverseIn[31];
  assign count[0] = \Bit_29_.countSoFar_0  | oneLeastReverseIn[31];

endmodule



module iNToRawFN_intWidth32
(
  signedIn,
  in,
  isZero,
  sign,
  sExp,
  sig
);

  input [31:0] in;
  output [7:0] sExp;
  output [32:0] sig;
  input signedIn;
  output isZero;
  output sign;
  wire [7:0] sExp;
  wire [32:0] sig;
  wire isZero,sign,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34;
  wire [31:0] absIn;
  wire [4:0] adjustedNormDist;
  assign sExp[6] = 1'b1;
  assign sExp[5] = 1'b0;
  assign sExp[7] = 1'b0;

  countLeadingZeros_inWidth32_countWidth5
  countLeadingZeros
  (
    .in(absIn),
    .count(adjustedNormDist)
  );

  assign sig = { 1'b0, absIn } << adjustedNormDist;
  assign { N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } = 1'b0 - in;
  assign absIn = (N0)? { N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } : 
                 (N1)? in : 1'b0;
  assign N0 = sign;
  assign N1 = N2;
  assign sign = signedIn & in[31];
  assign N2 = ~sign;
  assign isZero = ~sig[31];
  assign sExp[4] = ~adjustedNormDist[4];
  assign sExp[3] = ~adjustedNormDist[3];
  assign sExp[2] = ~adjustedNormDist[2];
  assign sExp[1] = ~adjustedNormDist[1];
  assign sExp[0] = ~adjustedNormDist[0];

endmodule



module roundAnyRawFNToRecFN_inExpWidth6_inSigWidth32_outExpWidth8_outSigWidth24_options5
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [7:0] in_sExp;
  input [32:0] in_sig;
  input [2:0] roundingMode;
  output [32:0] out;
  output [4:0] exceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [32:0] out;
  wire [4:0] exceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,exceptionFlags_4_,exceptionFlags_3_,roundMagUp,
  isNaNOut,\genblk2.roundPosBit ,\genblk2.anyRoundExtra ,\genblk2.anyRound ,
  \genblk2.roundIncr ,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,
  N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,
  N137,N138,N139,N140,common_inexact,notNaN_isSpecialInfOut,commonCase,
  overflow_roundMagUp,pegMinNonzeroMagOut,pegMaxFiniteMagOut,notNaN_isInfOut,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368;
  wire [8:0] sAdjustedExp,\genblk2.sRoundedExp ;
  wire [0:0] adjustedSig;
  wire [26:0] \genblk2.roundPosMask ;
  wire [25:0] \genblk2.roundedSig ;
  wire [22:0] common_fractOut;
  assign exceptionFlags_4_ = invalidExc;
  assign exceptionFlags[4] = exceptionFlags_4_;
  assign exceptionFlags_3_ = infiniteExc;
  assign exceptionFlags[3] = exceptionFlags_3_;
  assign N169 = ~roundingMode[2];
  assign N170 = roundingMode[1] | N169;
  assign N171 = roundingMode[0] | N170;
  assign N172 = ~N171;
  assign N173 = roundingMode[1] | roundingMode[2];
  assign N174 = roundingMode[0] | N173;
  assign N175 = ~N174;
  assign N176 = ~roundingMode[1];
  assign N177 = N176 | N169;
  assign N178 = roundingMode[0] | N177;
  assign N179 = ~N178;
  assign N180 = N176 | roundingMode[2];
  assign N181 = roundingMode[0] | N180;
  assign N182 = ~N181;
  assign N183 = ~roundingMode[0];
  assign N184 = N183 | N180;
  assign N185 = ~N184;
  assign sAdjustedExp = $signed(in_sExp) + $signed({ 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 });
  assign { N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36 } = { N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35 } + 1'b1;
  assign \genblk2.sRoundedExp  = sAdjustedExp + \genblk2.roundedSig [25:24];
  assign { N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90 } = (N0)? \genblk2.roundPosMask [26:1] : 
                                                                                                                                                                (N89)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N88;
  assign \genblk2.roundedSig  = (N1)? { N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87 } : 
                                (N2)? { N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140 } : 1'b0;
  assign N1 = \genblk2.roundIncr ;
  assign N2 = N9;
  assign common_fractOut = (N3)? \genblk2.roundedSig [23:1] : 
                           (N4)? \genblk2.roundedSig [22:0] : 1'b0;
  assign N3 = 1'b0;
  assign N4 = N196;
  assign out[32] = (N5)? 1'b0 : 
                   (N6)? in_sign : 1'b0;
  assign N5 = isNaNOut;
  assign N6 = N335;
  assign N144 = (N7)? common_fractOut[22] : 
                (N143)? 1'b0 : 1'b0;
  assign N7 = N142;
  assign { N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147 } = (N8)? common_fractOut[21:0] : 
                                                                                                                                                  (N146)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N145;
  assign roundMagUp = N186 | N188;
  assign N186 = N182 & in_sign;
  assign N188 = N185 & N187;
  assign N187 = ~in_sign;
  assign isNaNOut = exceptionFlags_4_ | N190;
  assign N190 = N189 & in_isNaN;
  assign N189 = ~exceptionFlags_3_;
  assign adjustedSig[0] = N195 | in_sig[0];
  assign N195 = N194 | in_sig[1];
  assign N194 = N193 | in_sig[2];
  assign N193 = N192 | in_sig[3];
  assign N192 = N191 | in_sig[4];
  assign N191 = in_sig[6] | in_sig[5];
  assign \genblk2.roundPosMask [26] = N196 & 1'b0;
  assign N196 = ~1'b0;
  assign \genblk2.roundPosMask [25] = N196 & 1'b0;
  assign \genblk2.roundPosMask [24] = N196 & 1'b0;
  assign \genblk2.roundPosMask [23] = N196 & 1'b0;
  assign \genblk2.roundPosMask [22] = N196 & 1'b0;
  assign \genblk2.roundPosMask [21] = N196 & 1'b0;
  assign \genblk2.roundPosMask [20] = N196 & 1'b0;
  assign \genblk2.roundPosMask [19] = N196 & 1'b0;
  assign \genblk2.roundPosMask [18] = N196 & 1'b0;
  assign \genblk2.roundPosMask [17] = N196 & 1'b0;
  assign \genblk2.roundPosMask [16] = N196 & 1'b0;
  assign \genblk2.roundPosMask [15] = N196 & 1'b0;
  assign \genblk2.roundPosMask [14] = N196 & 1'b0;
  assign \genblk2.roundPosMask [13] = N196 & 1'b0;
  assign \genblk2.roundPosMask [12] = N196 & 1'b0;
  assign \genblk2.roundPosMask [11] = N196 & 1'b0;
  assign \genblk2.roundPosMask [10] = N196 & 1'b0;
  assign \genblk2.roundPosMask [9] = N196 & 1'b0;
  assign \genblk2.roundPosMask [8] = N196 & 1'b0;
  assign \genblk2.roundPosMask [7] = N196 & 1'b0;
  assign \genblk2.roundPosMask [6] = N196 & 1'b0;
  assign \genblk2.roundPosMask [5] = N196 & 1'b0;
  assign \genblk2.roundPosMask [4] = N196 & 1'b0;
  assign \genblk2.roundPosMask [3] = N196 & 1'b0;
  assign \genblk2.roundPosMask [2] = N196 & 1'b0;
  assign \genblk2.roundPosMask [1] = N196 & 1'b1;
  assign \genblk2.roundPosMask [0] = N197 & 1'b1;
  assign N197 = ~1'b1;
  assign \genblk2.roundPosBit  = N244 | N250;
  assign N244 = N242 | N243;
  assign N242 = N240 | N241;
  assign N240 = N238 | N239;
  assign N238 = N236 | N237;
  assign N236 = N234 | N235;
  assign N234 = N232 | N233;
  assign N232 = N230 | N231;
  assign N230 = N228 | N229;
  assign N228 = N226 | N227;
  assign N226 = N224 | N225;
  assign N224 = N222 | N223;
  assign N222 = N220 | N221;
  assign N220 = N218 | N219;
  assign N218 = N216 | N217;
  assign N216 = N214 | N215;
  assign N214 = N212 | N213;
  assign N212 = N210 | N211;
  assign N210 = N208 | N209;
  assign N208 = N206 | N207;
  assign N206 = N204 | N205;
  assign N204 = N202 | N203;
  assign N202 = N200 | N201;
  assign N200 = N198 | N199;
  assign N198 = in_sig[32] & \genblk2.roundPosMask [26];
  assign N199 = in_sig[31] & \genblk2.roundPosMask [25];
  assign N201 = in_sig[30] & \genblk2.roundPosMask [24];
  assign N203 = in_sig[29] & \genblk2.roundPosMask [23];
  assign N205 = in_sig[28] & \genblk2.roundPosMask [22];
  assign N207 = in_sig[27] & \genblk2.roundPosMask [21];
  assign N209 = in_sig[26] & \genblk2.roundPosMask [20];
  assign N211 = in_sig[25] & \genblk2.roundPosMask [19];
  assign N213 = in_sig[24] & \genblk2.roundPosMask [18];
  assign N215 = in_sig[23] & \genblk2.roundPosMask [17];
  assign N217 = in_sig[22] & \genblk2.roundPosMask [16];
  assign N219 = in_sig[21] & \genblk2.roundPosMask [15];
  assign N221 = in_sig[20] & \genblk2.roundPosMask [14];
  assign N223 = in_sig[19] & \genblk2.roundPosMask [13];
  assign N225 = in_sig[18] & \genblk2.roundPosMask [12];
  assign N227 = in_sig[17] & \genblk2.roundPosMask [11];
  assign N229 = in_sig[16] & \genblk2.roundPosMask [10];
  assign N231 = in_sig[15] & \genblk2.roundPosMask [9];
  assign N233 = in_sig[14] & \genblk2.roundPosMask [8];
  assign N235 = in_sig[13] & \genblk2.roundPosMask [7];
  assign N237 = in_sig[12] & \genblk2.roundPosMask [6];
  assign N239 = in_sig[11] & \genblk2.roundPosMask [5];
  assign N241 = in_sig[10] & \genblk2.roundPosMask [4];
  assign N243 = in_sig[9] & \genblk2.roundPosMask [3];
  assign N250 = N249 & N196;
  assign N249 = N247 | N248;
  assign N247 = N245 | N246;
  assign N245 = in_sig[8] & \genblk2.roundPosMask [2];
  assign N246 = in_sig[7] & \genblk2.roundPosMask [1];
  assign N248 = adjustedSig[0] & \genblk2.roundPosMask [0];
  assign \genblk2.anyRoundExtra  = N297 | N303;
  assign N297 = N295 | N296;
  assign N295 = N293 | N294;
  assign N293 = N291 | N292;
  assign N291 = N289 | N290;
  assign N289 = N287 | N288;
  assign N287 = N285 | N286;
  assign N285 = N283 | N284;
  assign N283 = N281 | N282;
  assign N281 = N279 | N280;
  assign N279 = N277 | N278;
  assign N277 = N275 | N276;
  assign N275 = N273 | N274;
  assign N273 = N271 | N272;
  assign N271 = N269 | N270;
  assign N269 = N267 | N268;
  assign N267 = N265 | N266;
  assign N265 = N263 | N264;
  assign N263 = N261 | N262;
  assign N261 = N259 | N260;
  assign N259 = N257 | N258;
  assign N257 = N255 | N256;
  assign N255 = N253 | N254;
  assign N253 = N251 | N252;
  assign N251 = in_sig[32] & 1'b0;
  assign N252 = in_sig[31] & 1'b0;
  assign N254 = in_sig[30] & 1'b0;
  assign N256 = in_sig[29] & 1'b0;
  assign N258 = in_sig[28] & 1'b0;
  assign N260 = in_sig[27] & 1'b0;
  assign N262 = in_sig[26] & 1'b0;
  assign N264 = in_sig[25] & 1'b0;
  assign N266 = in_sig[24] & 1'b0;
  assign N268 = in_sig[23] & 1'b0;
  assign N270 = in_sig[22] & 1'b0;
  assign N272 = in_sig[21] & 1'b0;
  assign N274 = in_sig[20] & 1'b0;
  assign N276 = in_sig[19] & 1'b0;
  assign N278 = in_sig[18] & 1'b0;
  assign N280 = in_sig[17] & 1'b0;
  assign N282 = in_sig[16] & 1'b0;
  assign N284 = in_sig[15] & 1'b0;
  assign N286 = in_sig[14] & 1'b0;
  assign N288 = in_sig[13] & 1'b0;
  assign N290 = in_sig[12] & 1'b0;
  assign N292 = in_sig[11] & 1'b0;
  assign N294 = in_sig[10] & 1'b0;
  assign N296 = in_sig[9] & 1'b0;
  assign N303 = N302 & N196;
  assign N302 = N300 | N301;
  assign N300 = N298 | N299;
  assign N298 = in_sig[8] & 1'b0;
  assign N299 = in_sig[7] & 1'b0;
  assign N301 = adjustedSig[0] & 1'b1;
  assign \genblk2.anyRound  = \genblk2.roundPosBit  | \genblk2.anyRoundExtra ;
  assign \genblk2.roundIncr  = N305 | N306;
  assign N305 = N304 & \genblk2.roundPosBit ;
  assign N304 = N175 | N172;
  assign N306 = roundMagUp & \genblk2.anyRound ;
  assign N9 = ~\genblk2.roundIncr ;
  assign N10 = N307 & N308;
  assign N307 = N175 & \genblk2.roundPosBit ;
  assign N308 = ~\genblk2.anyRoundExtra ;
  assign N11 = in_sig[32] | 1'b0;
  assign N12 = in_sig[31] | 1'b0;
  assign N13 = in_sig[30] | 1'b0;
  assign N14 = in_sig[29] | 1'b0;
  assign N15 = in_sig[28] | 1'b0;
  assign N16 = in_sig[27] | 1'b0;
  assign N17 = in_sig[26] | 1'b0;
  assign N18 = in_sig[25] | 1'b0;
  assign N19 = in_sig[24] | 1'b0;
  assign N20 = in_sig[23] | 1'b0;
  assign N21 = in_sig[22] | 1'b0;
  assign N22 = in_sig[21] | 1'b0;
  assign N23 = in_sig[20] | 1'b0;
  assign N24 = in_sig[19] | 1'b0;
  assign N25 = in_sig[18] | 1'b0;
  assign N26 = in_sig[17] | 1'b0;
  assign N27 = in_sig[16] | 1'b0;
  assign N28 = in_sig[15] | 1'b0;
  assign N29 = in_sig[14] | 1'b0;
  assign N30 = in_sig[13] | 1'b0;
  assign N31 = in_sig[12] | 1'b0;
  assign N32 = in_sig[11] | 1'b0;
  assign N33 = in_sig[10] | 1'b0;
  assign N34 = in_sig[9] | 1'b0;
  assign N35 = in_sig[8] | 1'b0;
  assign N62 = N61 & N196;
  assign N63 = N60 & N196;
  assign N64 = N59 & N196;
  assign N65 = N58 & N196;
  assign N66 = N57 & N196;
  assign N67 = N56 & N196;
  assign N68 = N55 & N196;
  assign N69 = N54 & N196;
  assign N70 = N53 & N196;
  assign N71 = N52 & N196;
  assign N72 = N51 & N196;
  assign N73 = N50 & N196;
  assign N74 = N49 & N196;
  assign N75 = N48 & N196;
  assign N76 = N47 & N196;
  assign N77 = N46 & N196;
  assign N78 = N45 & N196;
  assign N79 = N44 & N196;
  assign N80 = N43 & N196;
  assign N81 = N42 & N196;
  assign N82 = N41 & N196;
  assign N83 = N40 & N196;
  assign N84 = N39 & N196;
  assign N85 = N38 & N196;
  assign N86 = N37 & N196;
  assign N87 = N36 & N309;
  assign N309 = ~N10;
  assign N88 = N179 & \genblk2.anyRound ;
  assign N89 = ~N88;
  assign N116 = N310 | N114;
  assign N310 = in_sig[32] & N196;
  assign N117 = N311 | N113;
  assign N311 = in_sig[31] & N196;
  assign N118 = N312 | N112;
  assign N312 = in_sig[30] & N196;
  assign N119 = N313 | N111;
  assign N313 = in_sig[29] & N196;
  assign N120 = N314 | N110;
  assign N314 = in_sig[28] & N196;
  assign N121 = N315 | N109;
  assign N315 = in_sig[27] & N196;
  assign N122 = N316 | N108;
  assign N316 = in_sig[26] & N196;
  assign N123 = N317 | N107;
  assign N317 = in_sig[25] & N196;
  assign N124 = N318 | N106;
  assign N318 = in_sig[24] & N196;
  assign N125 = N319 | N105;
  assign N319 = in_sig[23] & N196;
  assign N126 = N320 | N104;
  assign N320 = in_sig[22] & N196;
  assign N127 = N321 | N103;
  assign N321 = in_sig[21] & N196;
  assign N128 = N322 | N102;
  assign N322 = in_sig[20] & N196;
  assign N129 = N323 | N101;
  assign N323 = in_sig[19] & N196;
  assign N130 = N324 | N100;
  assign N324 = in_sig[18] & N196;
  assign N131 = N325 | N99;
  assign N325 = in_sig[17] & N196;
  assign N132 = N326 | N98;
  assign N326 = in_sig[16] & N196;
  assign N133 = N327 | N97;
  assign N327 = in_sig[15] & N196;
  assign N134 = N328 | N96;
  assign N328 = in_sig[14] & N196;
  assign N135 = N329 | N95;
  assign N329 = in_sig[13] & N196;
  assign N136 = N330 | N94;
  assign N330 = in_sig[12] & N196;
  assign N137 = N331 | N93;
  assign N331 = in_sig[11] & N196;
  assign N138 = N332 | N92;
  assign N332 = in_sig[10] & N196;
  assign N139 = N333 | N91;
  assign N333 = in_sig[9] & N196;
  assign N140 = N334 | N90;
  assign N334 = in_sig[8] & N196;
  assign common_inexact = 1'b0 | \genblk2.anyRound ;
  assign notNaN_isSpecialInfOut = exceptionFlags_3_ | in_isInf;
  assign commonCase = N337 & N338;
  assign N337 = N335 & N336;
  assign N335 = ~isNaNOut;
  assign N336 = ~notNaN_isSpecialInfOut;
  assign N338 = ~in_isZero;
  assign exceptionFlags[2] = commonCase & 1'b0;
  assign exceptionFlags[1] = commonCase & 1'b0;
  assign exceptionFlags[0] = exceptionFlags[2] | N339;
  assign N339 = commonCase & common_inexact;
  assign overflow_roundMagUp = N340 | roundMagUp;
  assign N340 = N175 | N172;
  assign pegMinNonzeroMagOut = N341 & N342;
  assign N341 = commonCase & 1'b0;
  assign N342 = roundMagUp | N179;
  assign pegMaxFiniteMagOut = exceptionFlags[2] & N343;
  assign N343 = ~overflow_roundMagUp;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | N344;
  assign N344 = exceptionFlags[2] & overflow_roundMagUp;
  assign N141 = in_isZero | 1'b0;
  assign out[31] = N350 | isNaNOut;
  assign N350 = N349 | notNaN_isInfOut;
  assign N349 = N348 | pegMaxFiniteMagOut;
  assign N348 = N346 & N347;
  assign N346 = \genblk2.sRoundedExp [8] & N345;
  assign N345 = ~N141;
  assign N347 = ~pegMinNonzeroMagOut;
  assign out[30] = N355 | isNaNOut;
  assign N355 = N354 | notNaN_isInfOut;
  assign N354 = N352 & N353;
  assign N352 = N351 & N347;
  assign N351 = \genblk2.sRoundedExp [7] & N345;
  assign N353 = ~pegMaxFiniteMagOut;
  assign out[29] = N360 | isNaNOut;
  assign N360 = N359 | pegMaxFiniteMagOut;
  assign N359 = N358 | pegMinNonzeroMagOut;
  assign N358 = N356 & N357;
  assign N356 = \genblk2.sRoundedExp [6] & N345;
  assign N357 = ~notNaN_isInfOut;
  assign out[28] = N361 | pegMaxFiniteMagOut;
  assign N361 = \genblk2.sRoundedExp [5] | pegMinNonzeroMagOut;
  assign out[27] = N362 | pegMaxFiniteMagOut;
  assign N362 = \genblk2.sRoundedExp [4] & N347;
  assign out[26] = N363 | pegMaxFiniteMagOut;
  assign N363 = \genblk2.sRoundedExp [3] | pegMinNonzeroMagOut;
  assign out[25] = N364 | pegMaxFiniteMagOut;
  assign N364 = \genblk2.sRoundedExp [2] & N347;
  assign out[24] = N365 | pegMaxFiniteMagOut;
  assign N365 = \genblk2.sRoundedExp [1] | pegMinNonzeroMagOut;
  assign out[23] = N366 | pegMaxFiniteMagOut;
  assign N366 = \genblk2.sRoundedExp [0] | pegMinNonzeroMagOut;
  assign N142 = N338 & N196;
  assign N143 = ~N142;
  assign N145 = N367 & N196;
  assign N367 = N335 & N338;
  assign N146 = ~N145;
  assign out[22] = N368 | pegMaxFiniteMagOut;
  assign N368 = isNaNOut | N144;
  assign out[21] = N168 | pegMaxFiniteMagOut;
  assign out[20] = N167 | pegMaxFiniteMagOut;
  assign out[19] = N166 | pegMaxFiniteMagOut;
  assign out[18] = N165 | pegMaxFiniteMagOut;
  assign out[17] = N164 | pegMaxFiniteMagOut;
  assign out[16] = N163 | pegMaxFiniteMagOut;
  assign out[15] = N162 | pegMaxFiniteMagOut;
  assign out[14] = N161 | pegMaxFiniteMagOut;
  assign out[13] = N160 | pegMaxFiniteMagOut;
  assign out[12] = N159 | pegMaxFiniteMagOut;
  assign out[11] = N158 | pegMaxFiniteMagOut;
  assign out[10] = N157 | pegMaxFiniteMagOut;
  assign out[9] = N156 | pegMaxFiniteMagOut;
  assign out[8] = N155 | pegMaxFiniteMagOut;
  assign out[7] = N154 | pegMaxFiniteMagOut;
  assign out[6] = N153 | pegMaxFiniteMagOut;
  assign out[5] = N152 | pegMaxFiniteMagOut;
  assign out[4] = N151 | pegMaxFiniteMagOut;
  assign out[3] = N150 | pegMaxFiniteMagOut;
  assign out[2] = N149 | pegMaxFiniteMagOut;
  assign out[1] = N148 | pegMaxFiniteMagOut;
  assign out[0] = N147 | pegMaxFiniteMagOut;

endmodule



module iNToRecFN_intWidth32_expWidth8_sigWidth24
(
  control,
  signedIn,
  in,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [31:0] in;
  input [2:0] roundingMode;
  output [32:0] out;
  output [4:0] exceptionFlags;
  input signedIn;
  wire [32:0] out,sig;
  wire [4:0] exceptionFlags;
  wire isZero,sign;
  wire [7:0] sExp;

  iNToRawFN_intWidth32
  iNToRawFN
  (
    .signedIn(signedIn),
    .in(in),
    .isZero(isZero),
    .sign(sign),
    .sExp(sExp),
    .sig(sig)
  );


  roundAnyRawFNToRecFN_inExpWidth6_inSigWidth32_outExpWidth8_outSigWidth24_options5
  roundRawToOut
  (
    .control(control[0]),
    .invalidExc(1'b0),
    .infiniteExc(1'b0),
    .in_isNaN(1'b0),
    .in_isInf(1'b0),
    .in_isZero(isZero),
    .in_sign(sign),
    .in_sExp(sExp),
    .in_sig(sig),
    .roundingMode(roundingMode),
    .out(out),
    .exceptionFlags(exceptionFlags)
  );


endmodule



module compareRecFN_expWidth8_sigWidth24
(
  a,
  b,
  signaling,
  lt,
  eq,
  gt,
  unordered,
  exceptionFlags
);

  input [32:0] a;
  input [32:0] b;
  output [4:0] exceptionFlags;
  input signaling;
  output lt;
  output eq;
  output gt;
  output unordered;
  wire [4:0] exceptionFlags;
  wire lt,eq,gt,unordered,N0,isNaNA,isInfA,isZeroA,signA,isSigNaNA,isNaNB,isInfB,
  isZeroB,signB,isSigNaNB,ordered,bothInfs,bothZeros,eqHiExps,N1,eqExps,N2,N3,N4,
  common_ltMags,N5,common_eqMags,ordered_lt,N6,ordered_eq,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31;
  wire [9:0] sExpA,sExpB;
  wire [24:0] sigA,sigB;
  assign exceptionFlags[0] = 1'b0;
  assign exceptionFlags[1] = 1'b0;
  assign exceptionFlags[2] = 1'b0;
  assign exceptionFlags[3] = 1'b0;

  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN_a
  (
    .in(a),
    .isNaN(isNaNA),
    .isInf(isInfA),
    .isZero(isZeroA),
    .sign(signA),
    .sExp(sExpA),
    .sig(sigA)
  );


  isSigNaNRecFN_expWidth8_sigWidth24
  isSigNaN_a
  (
    .in(a),
    .isSigNaN(isSigNaNA)
  );


  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN_b
  (
    .in(b),
    .isNaN(isNaNB),
    .isInf(isInfB),
    .isZero(isZeroB),
    .sign(signB),
    .sExp(sExpB),
    .sig(sigB)
  );


  isSigNaNRecFN_expWidth8_sigWidth24
  isSigNaN_b
  (
    .in(b),
    .isSigNaN(isSigNaNB)
  );

  assign eqHiExps = $signed({ 1'b0, sExpA[9:6] }) == $signed({ 1'b0, sExpB[9:6] });
  assign N1 = sExpA[5:0] == sExpB[5:0];
  assign N2 = $signed({ 1'b0, sExpA[9:6] }) < $signed({ 1'b0, sExpB[9:6] });
  assign N3 = sExpA[5:0] < sExpB[5:0];
  assign N4 = sigA < sigB;
  assign N5 = sigA == sigB;
  assign N0 = signA ^ signB;
  assign N6 = ~N0;
  assign ordered = N7 & N8;
  assign N7 = ~isNaNA;
  assign N8 = ~isNaNB;
  assign bothInfs = isInfA & isInfB;
  assign bothZeros = isZeroA & isZeroB;
  assign eqExps = eqHiExps & N1;
  assign common_ltMags = N10 | N11;
  assign N10 = N2 | N9;
  assign N9 = eqHiExps & N3;
  assign N11 = eqExps & N4;
  assign common_eqMags = eqExps & N5;
  assign ordered_lt = N12 & N23;
  assign N12 = ~bothZeros;
  assign N23 = N14 | N22;
  assign N14 = signA & N13;
  assign N13 = ~signB;
  assign N22 = N15 & N21;
  assign N15 = ~bothInfs;
  assign N21 = N19 | N20;
  assign N19 = N17 & N18;
  assign N17 = signA & N16;
  assign N16 = ~common_ltMags;
  assign N18 = ~common_eqMags;
  assign N20 = N13 & common_ltMags;
  assign ordered_eq = bothZeros | N25;
  assign N25 = N6 & N24;
  assign N24 = bothInfs | common_eqMags;
  assign exceptionFlags[4] = N26 | N28;
  assign N26 = isSigNaNA | isSigNaNB;
  assign N28 = signaling & N27;
  assign N27 = ~ordered;
  assign lt = ordered & ordered_lt;
  assign eq = ordered & ordered_eq;
  assign gt = N30 & N31;
  assign N30 = ordered & N29;
  assign N29 = ~ordered_lt;
  assign N31 = ~ordered_eq;
  assign unordered = ~ordered;

endmodule



module fpu_fmin_fmax_exp_width_p8_sig_width_p24
(
  fp_rs1_i,
  fp_rs2_i,
  fmin_not_fmax_i,
  invalid_o,
  result_o
);

  input [32:0] fp_rs1_i;
  input [32:0] fp_rs2_i;
  output [32:0] result_o;
  input fmin_not_fmax_i;
  output invalid_o;
  wire [32:0] result_o;
  wire invalid_o,N0,N1,rs1_is_nan,rs2_is_nan,rs1_is_signan,rs2_is_signan,cmp_lt_lo,
  cmp_eq_lo,both_zero_diff_sign,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5;

  compareRecFN_expWidth8_sigWidth24
  cmp0
  (
    .a(fp_rs1_i),
    .b(fp_rs2_i),
    .signaling(1'b0),
    .lt(cmp_lt_lo),
    .eq(cmp_eq_lo),
    .exceptionFlags({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5 })
  );

  assign { N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13 } = (N0)? fp_rs2_i : 
                                                                                                                                                                                   (N12)? fp_rs1_i : 1'b0;
  assign N0 = N11;
  assign result_o = (N1)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                    (N47)? fp_rs2_i : 
                    (N50)? fp_rs1_i : 
                    (N53)? { N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13 } : 
                    (N56)? fp_rs2_i : 
                    (N10)? fp_rs1_i : 1'b0;
  assign N1 = N2;
  assign rs1_is_nan = N57 & fp_rs1_i[29];
  assign N57 = fp_rs1_i[31] & fp_rs1_i[30];
  assign rs2_is_nan = N58 & fp_rs2_i[29];
  assign N58 = fp_rs2_i[31] & fp_rs2_i[30];
  assign rs1_is_signan = rs1_is_nan & N59;
  assign N59 = ~fp_rs1_i[22];
  assign rs2_is_signan = rs2_is_nan & N60;
  assign N60 = ~fp_rs2_i[22];
  assign both_zero_diff_sign = cmp_eq_lo & N61;
  assign N61 = fp_rs1_i[32] ^ fp_rs2_i[32];
  assign N2 = rs1_is_nan & rs2_is_nan;
  assign N3 = rs1_is_nan & N62;
  assign N62 = ~rs2_is_nan;
  assign N4 = N63 & rs2_is_nan;
  assign N63 = ~rs1_is_nan;
  assign N5 = cmp_lt_lo ^ fmin_not_fmax_i;
  assign N6 = N3 | N2;
  assign N7 = N4 | N6;
  assign N8 = both_zero_diff_sign | N7;
  assign N9 = N5 | N8;
  assign N10 = ~N9;
  assign N11 = fmin_not_fmax_i ^ fp_rs1_i[32];
  assign N12 = ~N11;
  assign N46 = ~N2;
  assign N47 = N3 & N46;
  assign N48 = ~N3;
  assign N49 = N46 & N48;
  assign N50 = N4 & N49;
  assign N51 = ~N4;
  assign N52 = N49 & N51;
  assign N53 = both_zero_diff_sign & N52;
  assign N54 = ~both_zero_diff_sign;
  assign N55 = N52 & N54;
  assign N56 = N5 & N55;
  assign invalid_o = rs1_is_signan | rs2_is_signan;

endmodule



module reverse_width23
(
  in,
  out
);

  input [22:0] in;
  output [22:0] out;
  wire [22:0] out;
  assign out[22] = in[0];
  assign out[21] = in[1];
  assign out[20] = in[2];
  assign out[19] = in[3];
  assign out[18] = in[4];
  assign out[17] = in[5];
  assign out[16] = in[6];
  assign out[15] = in[7];
  assign out[14] = in[8];
  assign out[13] = in[9];
  assign out[12] = in[10];
  assign out[11] = in[11];
  assign out[10] = in[12];
  assign out[9] = in[13];
  assign out[8] = in[14];
  assign out[7] = in[15];
  assign out[6] = in[16];
  assign out[5] = in[17];
  assign out[4] = in[18];
  assign out[3] = in[19];
  assign out[2] = in[20];
  assign out[1] = in[21];
  assign out[0] = in[22];

endmodule



module countLeadingZeros_inWidth23_countWidth5
(
  in,
  count
);

  input [22:0] in;
  output [4:0] count;
  wire [4:0] count;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,\Bit_5_.countSoFar_0 ,\Bit_9_.countSoFar_0 ,\Bit_10_.countSoFar_1 ,
  \Bit_11_.countSoFar_3 ,\Bit_13_.countSoFar_0 ,\Bit_17_.countSoFar_0 ,
  \Bit_18_.countSoFar_1 ,\Bit_19_.countSoFar_4 ,\Bit_20_.countSoFar_2 ,\Bit_21_.countSoFar_2 ,
  \Bit_21_.countSoFar_0 ,\Bit_22_.countSoFar_4 ,sv2v_dc_1;
  wire [22:0] reverseIn;
  wire [23:1] oneLeastReverseIn;
  wire [0:0] \Bit_1_.countSoFar ;
  wire [1:1] \Bit_2_.countSoFar ;
  wire [1:0] \Bit_3_.countSoFar ,\Bit_11_.countSoFar ,\Bit_19_.countSoFar ;
  wire [2:2] \Bit_4_.countSoFar ,\Bit_5_.countSoFar ;
  wire [2:1] \Bit_6_.countSoFar ,\Bit_22_.countSoFar ;
  wire [2:0] \Bit_7_.countSoFar ,\Bit_15_.countSoFar ;
  wire [3:3] \Bit_8_.countSoFar ,\Bit_9_.countSoFar ,\Bit_10_.countSoFar ;
  wire [3:2] \Bit_12_.countSoFar ,\Bit_13_.countSoFar ;
  wire [3:1] \Bit_14_.countSoFar ;
  wire [4:4] \Bit_16_.countSoFar ,\Bit_17_.countSoFar ,\Bit_18_.countSoFar ,
  \Bit_20_.countSoFar ,\Bit_21_.countSoFar ;

  reverse_width23
  reverse_in
  (
    .in(in),
    .out(reverseIn)
  );

  assign { oneLeastReverseIn[23:23], N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, sv2v_dc_1 } = { N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22 } + 1'b1;
  assign N0 = ~reverseIn[22];
  assign N1 = ~reverseIn[21];
  assign N2 = ~reverseIn[20];
  assign N3 = ~reverseIn[19];
  assign N4 = ~reverseIn[18];
  assign N5 = ~reverseIn[17];
  assign N6 = ~reverseIn[16];
  assign N7 = ~reverseIn[15];
  assign N8 = ~reverseIn[14];
  assign N9 = ~reverseIn[13];
  assign N10 = ~reverseIn[12];
  assign N11 = ~reverseIn[11];
  assign N12 = ~reverseIn[10];
  assign N13 = ~reverseIn[9];
  assign N14 = ~reverseIn[8];
  assign N15 = ~reverseIn[7];
  assign N16 = ~reverseIn[6];
  assign N17 = ~reverseIn[5];
  assign N18 = ~reverseIn[4];
  assign N19 = ~reverseIn[3];
  assign N20 = ~reverseIn[2];
  assign N21 = ~reverseIn[1];
  assign N22 = ~reverseIn[0];
  assign oneLeastReverseIn[22] = reverseIn[22] & N44;
  assign oneLeastReverseIn[21] = reverseIn[21] & N43;
  assign oneLeastReverseIn[20] = reverseIn[20] & N42;
  assign oneLeastReverseIn[19] = reverseIn[19] & N41;
  assign oneLeastReverseIn[18] = reverseIn[18] & N40;
  assign oneLeastReverseIn[17] = reverseIn[17] & N39;
  assign oneLeastReverseIn[16] = reverseIn[16] & N38;
  assign oneLeastReverseIn[15] = reverseIn[15] & N37;
  assign oneLeastReverseIn[14] = reverseIn[14] & N36;
  assign oneLeastReverseIn[13] = reverseIn[13] & N35;
  assign oneLeastReverseIn[12] = reverseIn[12] & N34;
  assign oneLeastReverseIn[11] = reverseIn[11] & N33;
  assign oneLeastReverseIn[10] = reverseIn[10] & N32;
  assign oneLeastReverseIn[9] = reverseIn[9] & N31;
  assign oneLeastReverseIn[8] = reverseIn[8] & N30;
  assign oneLeastReverseIn[7] = reverseIn[7] & N29;
  assign oneLeastReverseIn[6] = reverseIn[6] & N28;
  assign oneLeastReverseIn[5] = reverseIn[5] & N27;
  assign oneLeastReverseIn[4] = reverseIn[4] & N26;
  assign oneLeastReverseIn[3] = reverseIn[3] & N25;
  assign oneLeastReverseIn[2] = reverseIn[2] & N24;
  assign oneLeastReverseIn[1] = reverseIn[1] & N23;
  assign \Bit_1_.countSoFar [0] = 1'b0 | oneLeastReverseIn[1];
  assign \Bit_2_.countSoFar [1] = 1'b0 | oneLeastReverseIn[2];
  assign \Bit_3_.countSoFar [1] = \Bit_2_.countSoFar [1] | oneLeastReverseIn[3];
  assign \Bit_3_.countSoFar [0] = \Bit_1_.countSoFar [0] | oneLeastReverseIn[3];
  assign \Bit_4_.countSoFar [2] = 1'b0 | oneLeastReverseIn[4];
  assign \Bit_5_.countSoFar [2] = \Bit_4_.countSoFar [2] | oneLeastReverseIn[5];
  assign \Bit_5_.countSoFar_0  = \Bit_3_.countSoFar [0] | oneLeastReverseIn[5];
  assign \Bit_6_.countSoFar [2] = \Bit_5_.countSoFar [2] | oneLeastReverseIn[6];
  assign \Bit_6_.countSoFar [1] = \Bit_3_.countSoFar [1] | oneLeastReverseIn[6];
  assign \Bit_7_.countSoFar [2] = \Bit_6_.countSoFar [2] | oneLeastReverseIn[7];
  assign \Bit_7_.countSoFar [1] = \Bit_6_.countSoFar [1] | oneLeastReverseIn[7];
  assign \Bit_7_.countSoFar [0] = \Bit_5_.countSoFar_0  | oneLeastReverseIn[7];
  assign \Bit_8_.countSoFar [3] = 1'b0 | oneLeastReverseIn[8];
  assign \Bit_9_.countSoFar [3] = \Bit_8_.countSoFar [3] | oneLeastReverseIn[9];
  assign \Bit_9_.countSoFar_0  = \Bit_7_.countSoFar [0] | oneLeastReverseIn[9];
  assign \Bit_10_.countSoFar [3] = \Bit_9_.countSoFar [3] | oneLeastReverseIn[10];
  assign \Bit_10_.countSoFar_1  = \Bit_7_.countSoFar [1] | oneLeastReverseIn[10];
  assign \Bit_11_.countSoFar_3  = \Bit_10_.countSoFar [3] | oneLeastReverseIn[11];
  assign \Bit_11_.countSoFar [1] = \Bit_10_.countSoFar_1  | oneLeastReverseIn[11];
  assign \Bit_11_.countSoFar [0] = \Bit_9_.countSoFar_0  | oneLeastReverseIn[11];
  assign \Bit_12_.countSoFar [3] = \Bit_11_.countSoFar_3  | oneLeastReverseIn[12];
  assign \Bit_12_.countSoFar [2] = \Bit_7_.countSoFar [2] | oneLeastReverseIn[12];
  assign \Bit_13_.countSoFar [3] = \Bit_12_.countSoFar [3] | oneLeastReverseIn[13];
  assign \Bit_13_.countSoFar [2] = \Bit_12_.countSoFar [2] | oneLeastReverseIn[13];
  assign \Bit_13_.countSoFar_0  = \Bit_11_.countSoFar [0] | oneLeastReverseIn[13];
  assign \Bit_14_.countSoFar [3] = \Bit_13_.countSoFar [3] | oneLeastReverseIn[14];
  assign \Bit_14_.countSoFar [2] = \Bit_13_.countSoFar [2] | oneLeastReverseIn[14];
  assign \Bit_14_.countSoFar [1] = \Bit_11_.countSoFar [1] | oneLeastReverseIn[14];
  assign count[3] = \Bit_14_.countSoFar [3] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [2] = \Bit_14_.countSoFar [2] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [1] = \Bit_14_.countSoFar [1] | oneLeastReverseIn[15];
  assign \Bit_15_.countSoFar [0] = \Bit_13_.countSoFar_0  | oneLeastReverseIn[15];
  assign \Bit_16_.countSoFar [4] = 1'b0 | oneLeastReverseIn[16];
  assign \Bit_17_.countSoFar [4] = \Bit_16_.countSoFar [4] | oneLeastReverseIn[17];
  assign \Bit_17_.countSoFar_0  = \Bit_15_.countSoFar [0] | oneLeastReverseIn[17];
  assign \Bit_18_.countSoFar [4] = \Bit_17_.countSoFar [4] | oneLeastReverseIn[18];
  assign \Bit_18_.countSoFar_1  = \Bit_15_.countSoFar [1] | oneLeastReverseIn[18];
  assign \Bit_19_.countSoFar_4  = \Bit_18_.countSoFar [4] | oneLeastReverseIn[19];
  assign \Bit_19_.countSoFar [1] = \Bit_18_.countSoFar_1  | oneLeastReverseIn[19];
  assign \Bit_19_.countSoFar [0] = \Bit_17_.countSoFar_0  | oneLeastReverseIn[19];
  assign \Bit_20_.countSoFar [4] = \Bit_19_.countSoFar_4  | oneLeastReverseIn[20];
  assign \Bit_20_.countSoFar_2  = \Bit_15_.countSoFar [2] | oneLeastReverseIn[20];
  assign \Bit_21_.countSoFar [4] = \Bit_20_.countSoFar [4] | oneLeastReverseIn[21];
  assign \Bit_21_.countSoFar_2  = \Bit_20_.countSoFar_2  | oneLeastReverseIn[21];
  assign \Bit_21_.countSoFar_0  = \Bit_19_.countSoFar [0] | oneLeastReverseIn[21];
  assign \Bit_22_.countSoFar_4  = \Bit_21_.countSoFar [4] | oneLeastReverseIn[22];
  assign \Bit_22_.countSoFar [2] = \Bit_21_.countSoFar_2  | oneLeastReverseIn[22];
  assign \Bit_22_.countSoFar [1] = \Bit_19_.countSoFar [1] | oneLeastReverseIn[22];
  assign count[4] = \Bit_22_.countSoFar_4  | oneLeastReverseIn[23];
  assign count[2] = \Bit_22_.countSoFar [2] | oneLeastReverseIn[23];
  assign count[1] = \Bit_22_.countSoFar [1] | oneLeastReverseIn[23];
  assign count[0] = \Bit_21_.countSoFar_0  | oneLeastReverseIn[23];

endmodule



module fNToRecFN_expWidth8_sigWidth24
(
  in,
  out
);

  input [31:0] in;
  output [32:0] out;
  wire [32:0] out;
  wire N0,N1,N2,out_32_,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,isZero,isSpecial,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50;
  wire [4:0] normDist;
  wire [22:1] subnormFract;
  wire [8:6] adjustedExp;
  assign out_32_ = in[31];
  assign out[32] = out_32_;

  countLeadingZeros_inWidth23_countWidth5
  countLeadingZeros
  (
    .in(in[22:0]),
    .count(normDist)
  );

  assign isSpecial = adjustedExp[8:7] == { 1'b1, 1'b1 };
  assign subnormFract = in[21:0] << normDist;
  assign N20 = in[21] | in[22];
  assign N21 = in[20] | N20;
  assign N22 = in[19] | N21;
  assign N23 = in[18] | N22;
  assign N24 = in[17] | N23;
  assign N25 = in[16] | N24;
  assign N26 = in[15] | N25;
  assign N27 = in[14] | N26;
  assign N28 = in[13] | N27;
  assign N29 = in[12] | N28;
  assign N30 = in[11] | N29;
  assign N31 = in[10] | N30;
  assign N32 = in[9] | N31;
  assign N33 = in[8] | N32;
  assign N34 = in[7] | N33;
  assign N35 = in[6] | N34;
  assign N36 = in[5] | N35;
  assign N37 = in[4] | N36;
  assign N38 = in[3] | N37;
  assign N39 = in[2] | N38;
  assign N40 = in[1] | N39;
  assign N41 = in[0] | N40;
  assign N42 = ~N41;
  assign N43 = in[29] | in[30];
  assign N44 = in[28] | N43;
  assign N45 = in[27] | N44;
  assign N46 = in[26] | N45;
  assign N47 = in[25] | N46;
  assign N48 = in[24] | N47;
  assign N49 = in[23] | N48;
  assign N50 = ~N49;
  assign { adjustedExp, out[28:23] } = { N50, N15, N14, N13, N12, N11, N10, N9, N8 } + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N50, N49 };
  assign { N15, N14, N13, N12, N11, N10, N9, N8 } = (N0)? { 1'b1, 1'b1, 1'b1, N3, N4, N5, N6, N7 } : 
                                                    (N1)? in[30:23] : 1'b0;
  assign N0 = N50;
  assign N1 = N49;
  assign out[31:29] = (N2)? { 1'b1, 1'b1, N41 } : 
                      (N19)? { 1'b0, 1'b0, 1'b0 } : 
                      (N17)? adjustedExp : 1'b0;
  assign N2 = isSpecial;
  assign out[22:0] = (N0)? { subnormFract, 1'b0 } : 
                     (N1)? in[22:0] : 1'b0;
  assign N3 = ~normDist[4];
  assign N4 = ~normDist[3];
  assign N5 = ~normDist[2];
  assign N6 = ~normDist[1];
  assign N7 = ~normDist[0];
  assign isZero = N50 & N42;
  assign N16 = isZero | isSpecial;
  assign N17 = ~N16;
  assign N18 = ~isSpecial;
  assign N19 = isZero & N18;

endmodule



module fpu_float_aux
(
  fp_v_i,
  fpu_float_op_i,
  fp_rs1_i,
  fp_rs2_i,
  fp_rm_i,
  v_o,
  result_o,
  fflags_o_invalid_,
  fflags_o_div_zero_,
  fflags_o_overflow_,
  fflags_o_underflow_,
  fflags_o_inexact_
);

  input [3:0] fpu_float_op_i;
  input [32:0] fp_rs1_i;
  input [32:0] fp_rs2_i;
  input [2:0] fp_rm_i;
  output [32:0] result_o;
  input fp_v_i;
  output v_o;
  output fflags_o_invalid_;
  output fflags_o_div_zero_;
  output fflags_o_overflow_;
  output fflags_o_underflow_;
  output fflags_o_inexact_;
  wire [32:0] result_o,i2f_result_lo,fmin_fmax_result_lo,rs1_recoded_val;
  wire v_o,fflags_o_invalid_,fflags_o_div_zero_,fflags_o_overflow_,fflags_o_underflow_,
  fflags_o_inexact_,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,i2f_fflags_lo_invalid_,
  i2f_fflags_lo_div_zero_,i2f_fflags_lo_overflow_,i2f_fflags_lo_underflow_,
  i2f_fflags_lo_inexact_,fmin_fmax_invalid_lo,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71;
  wire [32:32] fsgnj_result;

  iNToRecFN_intWidth32_expWidth8_sigWidth24
  i2f
  (
    .control(1'b1),
    .signedIn(N55),
    .in(fp_rs1_i[31:0]),
    .roundingMode(fp_rm_i),
    .out(i2f_result_lo),
    .exceptionFlags({ i2f_fflags_lo_invalid_, i2f_fflags_lo_div_zero_, i2f_fflags_lo_overflow_, i2f_fflags_lo_underflow_, i2f_fflags_lo_inexact_ })
  );


  fpu_fmin_fmax_exp_width_p8_sig_width_p24
  minmax0
  (
    .fp_rs1_i(fp_rs1_i),
    .fp_rs2_i(fp_rs2_i),
    .fmin_not_fmax_i(N61),
    .invalid_o(fmin_fmax_invalid_lo),
    .result_o(fmin_fmax_result_lo)
  );

  assign N10 = fpu_float_op_i[2] | N57;
  assign N11 = N10 | N48;
  assign N13 = N15 | fpu_float_op_i[0];
  assign N15 = N56 | fpu_float_op_i[1];
  assign N16 = N15 | N48;

  fNToRecFN_expWidth8_sigWidth24
  recFN_rs1
  (
    .in(fp_rs1_i[31:0]),
    .out(rs1_recoded_val)
  );

  assign N24 = fpu_float_op_i[3] | N56;
  assign N25 = N57 | fpu_float_op_i[0];
  assign N26 = N24 | N25;
  assign N27 = N57 | N48;
  assign N28 = N24 | N27;
  assign N30 = N51 | fpu_float_op_i[2];
  assign N31 = fpu_float_op_i[1] | fpu_float_op_i[0];
  assign N32 = N30 | N31;
  assign N33 = fpu_float_op_i[1] | N48;
  assign N34 = N30 | N33;
  assign N36 = fpu_float_op_i[3] | fpu_float_op_i[2];
  assign N37 = N36 | N27;
  assign N38 = N24 | N31;
  assign N39 = N24 | N33;
  assign N41 = N30 | N25;
  assign N43 = fpu_float_op_i[3] & fpu_float_op_i[1];
  assign N44 = N43 & fpu_float_op_i[0];
  assign N45 = N51 & N56;
  assign N46 = N45 & N57;
  assign N47 = fpu_float_op_i[3] & fpu_float_op_i[2];
  assign N49 = N45 & N48;
  assign N51 = ~fpu_float_op_i[3];
  assign N52 = fpu_float_op_i[2] | N51;
  assign N53 = fpu_float_op_i[1] | N52;
  assign N54 = fpu_float_op_i[0] | N53;
  assign N55 = ~N54;
  assign N56 = ~fpu_float_op_i[2];
  assign N57 = ~fpu_float_op_i[1];
  assign N58 = N56 | fpu_float_op_i[3];
  assign N59 = N57 | N58;
  assign N60 = fpu_float_op_i[0] | N59;
  assign N61 = ~N60;
  assign N23 = (N0)? fp_rs2_i[32] : 
               (N1)? N21 : 
               (N2)? N22 : 
               (N20)? fp_rs1_i[32] : 1'b0;
  assign N0 = N12;
  assign N1 = N14;
  assign N2 = N17;
  assign fsgnj_result[32] = (N3)? N23 : 
                            (N4)? fp_rs1_i[32] : 1'b0;
  assign N3 = N51;
  assign N4 = fpu_float_op_i[3];
  assign v_o = (N5)? fp_v_i : 
               (N6)? fp_v_i : 
               (N7)? fp_v_i : 
               (N8)? fp_v_i : 
               (N9)? 1'b0 : 1'b0;
  assign N5 = N29;
  assign N6 = N35;
  assign N7 = N40;
  assign N8 = N42;
  assign N9 = N50;
  assign result_o = (N5)? fmin_fmax_result_lo : 
                    (N6)? i2f_result_lo : 
                    (N7)? { fsgnj_result[32:32], fp_rs1_i[31:0] } : 
                    (N8)? rs1_recoded_val : 
                    (N9)? i2f_result_lo : 1'b0;
  assign { fflags_o_invalid_, fflags_o_div_zero_, fflags_o_overflow_, fflags_o_underflow_, fflags_o_inexact_ } = (N5)? { fmin_fmax_invalid_lo, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                 (N6)? { i2f_fflags_lo_invalid_, i2f_fflags_lo_div_zero_, i2f_fflags_lo_overflow_, i2f_fflags_lo_underflow_, i2f_fflags_lo_inexact_ } : 
                                                                                                                 (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                 (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                 (N9)? { i2f_fflags_lo_invalid_, i2f_fflags_lo_div_zero_, i2f_fflags_lo_overflow_, i2f_fflags_lo_underflow_, i2f_fflags_lo_inexact_ } : 1'b0;
  assign N12 = ~N11;
  assign N14 = ~N13;
  assign N17 = ~N16;
  assign N18 = N14 | N12;
  assign N19 = N17 | N18;
  assign N20 = ~N19;
  assign N21 = ~fp_rs2_i[32];
  assign N22 = fp_rs1_i[32] ^ fp_rs2_i[32];
  assign N29 = N62 | N63;
  assign N62 = ~N26;
  assign N63 = ~N28;
  assign N35 = N64 | N65;
  assign N64 = ~N32;
  assign N65 = ~N34;
  assign N40 = N68 | N69;
  assign N68 = N66 | N67;
  assign N66 = ~N37;
  assign N67 = ~N38;
  assign N69 = ~N39;
  assign N42 = ~N41;
  assign N48 = ~fpu_float_op_i[0];
  assign N50 = N44 | N71;
  assign N71 = N46 | N70;
  assign N70 = N47 | N49;

endmodule



module fpu_float
(
  clk_i,
  reset_i,
  stall_fpu1_i,
  stall_fpu2_i,
  imul_v_i,
  imul_rs1_i,
  imul_rs2_i,
  imul_rd_i,
  fp_v_i,
  fpu_float_op_i,
  fp_rs1_i,
  fp_rs2_i,
  fp_rs3_i,
  fp_rd_i,
  fp_rm_i,
  imul_v_o,
  imul_result_o,
  imul_rd_o,
  fp_v_o,
  fp_result_o,
  fp_rd_o,
  fpu1_v_r_o,
  fpu1_rd_o,
  fp_fflags_o_invalid_,
  fp_fflags_o_div_zero_,
  fp_fflags_o_overflow_,
  fp_fflags_o_underflow_,
  fp_fflags_o_inexact_
);

  input [31:0] imul_rs1_i;
  input [31:0] imul_rs2_i;
  input [4:0] imul_rd_i;
  input [3:0] fpu_float_op_i;
  input [32:0] fp_rs1_i;
  input [32:0] fp_rs2_i;
  input [32:0] fp_rs3_i;
  input [4:0] fp_rd_i;
  input [2:0] fp_rm_i;
  output [31:0] imul_result_o;
  output [4:0] imul_rd_o;
  output [32:0] fp_result_o;
  output [4:0] fp_rd_o;
  output [4:0] fpu1_rd_o;
  input clk_i;
  input reset_i;
  input stall_fpu1_i;
  input stall_fpu2_i;
  input imul_v_i;
  input fp_v_i;
  output imul_v_o;
  output fp_v_o;
  output fpu1_v_r_o;
  output fp_fflags_o_invalid_;
  output fp_fflags_o_div_zero_;
  output fp_fflags_o_overflow_;
  output fp_fflags_o_underflow_;
  output fp_fflags_o_inexact_;
  wire [31:0] imul_result_o;
  wire [4:0] imul_rd_o,fp_rd_o,fpu1_rd_o;
  wire [32:0] fp_result_o,fma2_result_lo,aux_result_lo;
  wire imul_v_o,fp_v_o,fpu1_v_r_o,fp_fflags_o_invalid_,fp_fflags_o_div_zero_,
  fp_fflags_o_overflow_,fp_fflags_o_underflow_,fp_fflags_o_inexact_,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,fma1_v_lo,invalidExc,out_isNaN,out_isInf,out_isZero,out_sign,
  fma2_v_lo,fma2_fflags_lo_invalid_,fma2_fflags_lo_div_zero_,fma2_fflags_lo_overflow_,
  fma2_fflags_lo_underflow_,fma2_fflags_lo_inexact_,aux_v_lo,aux_fflags_lo_invalid_,
  aux_fflags_lo_div_zero_,aux_fflags_lo_overflow_,aux_fflags_lo_underflow_,
  aux_fflags_lo_inexact_,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37;
  wire [2:0] fma1_rm_lo;
  wire [9:0] out_sExp,aux_fflags_r;
  wire [26:0] out_sig;
  wire [1:0] aux_v_r;
  wire [65:0] aux_result_r;
  reg fp_rd_o_4_sv2v_reg,fp_rd_o_3_sv2v_reg,fp_rd_o_2_sv2v_reg,fp_rd_o_1_sv2v_reg,
  fp_rd_o_0_sv2v_reg,fpu1_rd_o_4_sv2v_reg,fpu1_rd_o_3_sv2v_reg,fpu1_rd_o_2_sv2v_reg,
  fpu1_rd_o_1_sv2v_reg,fpu1_rd_o_0_sv2v_reg,aux_fflags_r_9_sv2v_reg,
  aux_fflags_r_8_sv2v_reg,aux_fflags_r_7_sv2v_reg,aux_fflags_r_6_sv2v_reg,aux_fflags_r_5_sv2v_reg,
  aux_fflags_r_4_sv2v_reg,aux_fflags_r_3_sv2v_reg,aux_fflags_r_2_sv2v_reg,
  aux_fflags_r_1_sv2v_reg,aux_fflags_r_0_sv2v_reg,aux_v_r_1_sv2v_reg,aux_v_r_0_sv2v_reg,
  aux_result_r_65_sv2v_reg,aux_result_r_64_sv2v_reg,aux_result_r_63_sv2v_reg,
  aux_result_r_62_sv2v_reg,aux_result_r_61_sv2v_reg,aux_result_r_60_sv2v_reg,
  aux_result_r_59_sv2v_reg,aux_result_r_58_sv2v_reg,aux_result_r_57_sv2v_reg,
  aux_result_r_56_sv2v_reg,aux_result_r_55_sv2v_reg,aux_result_r_54_sv2v_reg,
  aux_result_r_53_sv2v_reg,aux_result_r_52_sv2v_reg,aux_result_r_51_sv2v_reg,aux_result_r_50_sv2v_reg,
  aux_result_r_49_sv2v_reg,aux_result_r_48_sv2v_reg,aux_result_r_47_sv2v_reg,
  aux_result_r_46_sv2v_reg,aux_result_r_45_sv2v_reg,aux_result_r_44_sv2v_reg,
  aux_result_r_43_sv2v_reg,aux_result_r_42_sv2v_reg,aux_result_r_41_sv2v_reg,
  aux_result_r_40_sv2v_reg,aux_result_r_39_sv2v_reg,aux_result_r_38_sv2v_reg,
  aux_result_r_37_sv2v_reg,aux_result_r_36_sv2v_reg,aux_result_r_35_sv2v_reg,aux_result_r_34_sv2v_reg,
  aux_result_r_33_sv2v_reg,aux_result_r_32_sv2v_reg,aux_result_r_31_sv2v_reg,
  aux_result_r_30_sv2v_reg,aux_result_r_29_sv2v_reg,aux_result_r_28_sv2v_reg,
  aux_result_r_27_sv2v_reg,aux_result_r_26_sv2v_reg,aux_result_r_25_sv2v_reg,
  aux_result_r_24_sv2v_reg,aux_result_r_23_sv2v_reg,aux_result_r_22_sv2v_reg,
  aux_result_r_21_sv2v_reg,aux_result_r_20_sv2v_reg,aux_result_r_19_sv2v_reg,aux_result_r_18_sv2v_reg,
  aux_result_r_17_sv2v_reg,aux_result_r_16_sv2v_reg,aux_result_r_15_sv2v_reg,
  aux_result_r_14_sv2v_reg,aux_result_r_13_sv2v_reg,aux_result_r_12_sv2v_reg,
  aux_result_r_11_sv2v_reg,aux_result_r_10_sv2v_reg,aux_result_r_9_sv2v_reg,
  aux_result_r_8_sv2v_reg,aux_result_r_7_sv2v_reg,aux_result_r_6_sv2v_reg,aux_result_r_5_sv2v_reg,
  aux_result_r_4_sv2v_reg,aux_result_r_3_sv2v_reg,aux_result_r_2_sv2v_reg,
  aux_result_r_1_sv2v_reg,aux_result_r_0_sv2v_reg;
  assign fp_rd_o[4] = fp_rd_o_4_sv2v_reg;
  assign fp_rd_o[3] = fp_rd_o_3_sv2v_reg;
  assign fp_rd_o[2] = fp_rd_o_2_sv2v_reg;
  assign fp_rd_o[1] = fp_rd_o_1_sv2v_reg;
  assign fp_rd_o[0] = fp_rd_o_0_sv2v_reg;
  assign fpu1_rd_o[4] = fpu1_rd_o_4_sv2v_reg;
  assign fpu1_rd_o[3] = fpu1_rd_o_3_sv2v_reg;
  assign fpu1_rd_o[2] = fpu1_rd_o_2_sv2v_reg;
  assign fpu1_rd_o[1] = fpu1_rd_o_1_sv2v_reg;
  assign fpu1_rd_o[0] = fpu1_rd_o_0_sv2v_reg;
  assign aux_fflags_r[9] = aux_fflags_r_9_sv2v_reg;
  assign aux_fflags_r[8] = aux_fflags_r_8_sv2v_reg;
  assign aux_fflags_r[7] = aux_fflags_r_7_sv2v_reg;
  assign aux_fflags_r[6] = aux_fflags_r_6_sv2v_reg;
  assign aux_fflags_r[5] = aux_fflags_r_5_sv2v_reg;
  assign aux_fflags_r[4] = aux_fflags_r_4_sv2v_reg;
  assign aux_fflags_r[3] = aux_fflags_r_3_sv2v_reg;
  assign aux_fflags_r[2] = aux_fflags_r_2_sv2v_reg;
  assign aux_fflags_r[1] = aux_fflags_r_1_sv2v_reg;
  assign aux_fflags_r[0] = aux_fflags_r_0_sv2v_reg;
  assign aux_v_r[1] = aux_v_r_1_sv2v_reg;
  assign aux_v_r[0] = aux_v_r_0_sv2v_reg;
  assign aux_result_r[65] = aux_result_r_65_sv2v_reg;
  assign aux_result_r[64] = aux_result_r_64_sv2v_reg;
  assign aux_result_r[63] = aux_result_r_63_sv2v_reg;
  assign aux_result_r[62] = aux_result_r_62_sv2v_reg;
  assign aux_result_r[61] = aux_result_r_61_sv2v_reg;
  assign aux_result_r[60] = aux_result_r_60_sv2v_reg;
  assign aux_result_r[59] = aux_result_r_59_sv2v_reg;
  assign aux_result_r[58] = aux_result_r_58_sv2v_reg;
  assign aux_result_r[57] = aux_result_r_57_sv2v_reg;
  assign aux_result_r[56] = aux_result_r_56_sv2v_reg;
  assign aux_result_r[55] = aux_result_r_55_sv2v_reg;
  assign aux_result_r[54] = aux_result_r_54_sv2v_reg;
  assign aux_result_r[53] = aux_result_r_53_sv2v_reg;
  assign aux_result_r[52] = aux_result_r_52_sv2v_reg;
  assign aux_result_r[51] = aux_result_r_51_sv2v_reg;
  assign aux_result_r[50] = aux_result_r_50_sv2v_reg;
  assign aux_result_r[49] = aux_result_r_49_sv2v_reg;
  assign aux_result_r[48] = aux_result_r_48_sv2v_reg;
  assign aux_result_r[47] = aux_result_r_47_sv2v_reg;
  assign aux_result_r[46] = aux_result_r_46_sv2v_reg;
  assign aux_result_r[45] = aux_result_r_45_sv2v_reg;
  assign aux_result_r[44] = aux_result_r_44_sv2v_reg;
  assign aux_result_r[43] = aux_result_r_43_sv2v_reg;
  assign aux_result_r[42] = aux_result_r_42_sv2v_reg;
  assign aux_result_r[41] = aux_result_r_41_sv2v_reg;
  assign aux_result_r[40] = aux_result_r_40_sv2v_reg;
  assign aux_result_r[39] = aux_result_r_39_sv2v_reg;
  assign aux_result_r[38] = aux_result_r_38_sv2v_reg;
  assign aux_result_r[37] = aux_result_r_37_sv2v_reg;
  assign aux_result_r[36] = aux_result_r_36_sv2v_reg;
  assign aux_result_r[35] = aux_result_r_35_sv2v_reg;
  assign aux_result_r[34] = aux_result_r_34_sv2v_reg;
  assign aux_result_r[33] = aux_result_r_33_sv2v_reg;
  assign aux_result_r[32] = aux_result_r_32_sv2v_reg;
  assign aux_result_r[31] = aux_result_r_31_sv2v_reg;
  assign aux_result_r[30] = aux_result_r_30_sv2v_reg;
  assign aux_result_r[29] = aux_result_r_29_sv2v_reg;
  assign aux_result_r[28] = aux_result_r_28_sv2v_reg;
  assign aux_result_r[27] = aux_result_r_27_sv2v_reg;
  assign aux_result_r[26] = aux_result_r_26_sv2v_reg;
  assign aux_result_r[25] = aux_result_r_25_sv2v_reg;
  assign aux_result_r[24] = aux_result_r_24_sv2v_reg;
  assign aux_result_r[23] = aux_result_r_23_sv2v_reg;
  assign aux_result_r[22] = aux_result_r_22_sv2v_reg;
  assign aux_result_r[21] = aux_result_r_21_sv2v_reg;
  assign aux_result_r[20] = aux_result_r_20_sv2v_reg;
  assign aux_result_r[19] = aux_result_r_19_sv2v_reg;
  assign aux_result_r[18] = aux_result_r_18_sv2v_reg;
  assign aux_result_r[17] = aux_result_r_17_sv2v_reg;
  assign aux_result_r[16] = aux_result_r_16_sv2v_reg;
  assign aux_result_r[15] = aux_result_r_15_sv2v_reg;
  assign aux_result_r[14] = aux_result_r_14_sv2v_reg;
  assign aux_result_r[13] = aux_result_r_13_sv2v_reg;
  assign aux_result_r[12] = aux_result_r_12_sv2v_reg;
  assign aux_result_r[11] = aux_result_r_11_sv2v_reg;
  assign aux_result_r[10] = aux_result_r_10_sv2v_reg;
  assign aux_result_r[9] = aux_result_r_9_sv2v_reg;
  assign aux_result_r[8] = aux_result_r_8_sv2v_reg;
  assign aux_result_r[7] = aux_result_r_7_sv2v_reg;
  assign aux_result_r[6] = aux_result_r_6_sv2v_reg;
  assign aux_result_r[5] = aux_result_r_5_sv2v_reg;
  assign aux_result_r[4] = aux_result_r_4_sv2v_reg;
  assign aux_result_r[3] = aux_result_r_3_sv2v_reg;
  assign aux_result_r[2] = aux_result_r_2_sv2v_reg;
  assign aux_result_r[1] = aux_result_r_1_sv2v_reg;
  assign aux_result_r[0] = aux_result_r_0_sv2v_reg;
  assign imul_rd_o[4] = fpu1_rd_o[4];
  assign imul_rd_o[3] = fpu1_rd_o[3];
  assign imul_rd_o[2] = fpu1_rd_o[2];
  assign imul_rd_o[1] = fpu1_rd_o[1];
  assign imul_rd_o[0] = fpu1_rd_o[0];

  fpu_float_fma
  fma1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .stall_fpu1_i(stall_fpu1_i),
    .imul_v_i(imul_v_i),
    .imul_rs1_i(imul_rs1_i),
    .imul_rs2_i(imul_rs2_i),
    .fp_v_i(fp_v_i),
    .fpu_float_op_i(fpu_float_op_i),
    .fp_rs1_i(fp_rs1_i),
    .fp_rs2_i(fp_rs2_i),
    .fp_rs3_i(fp_rs3_i),
    .fp_rm_i(fp_rm_i),
    .imul_v_o(imul_v_o),
    .imul_result_o(imul_result_o),
    .fma1_v_o(fma1_v_lo),
    .fma1_rm_o(fma1_rm_lo),
    .invalidExc_o(invalidExc),
    .out_isNaN_o(out_isNaN),
    .out_isInf_o(out_isInf),
    .out_isZero_o(out_isZero),
    .out_sign_o(out_sign),
    .out_sExp_o(out_sExp),
    .out_sig_o(out_sig)
  );


  fpu_float_fma_round
  fma2
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .stall_fpu2_i(stall_fpu2_i),
    .fma1_v_i(fma1_v_lo),
    .fma1_rm_i(fma1_rm_lo),
    .invalidExc_i(invalidExc),
    .in_isNaN_i(out_isNaN),
    .in_isInf_i(out_isInf),
    .in_isZero_i(out_isZero),
    .in_sign_i(out_sign),
    .in_sExp_i(out_sExp),
    .in_sig_i(out_sig),
    .fma2_v_o(fma2_v_lo),
    .fma2_result_o(fma2_result_lo),
    .fma2_fflags_o_invalid_(fma2_fflags_lo_invalid_),
    .fma2_fflags_o_div_zero_(fma2_fflags_lo_div_zero_),
    .fma2_fflags_o_overflow_(fma2_fflags_lo_overflow_),
    .fma2_fflags_o_underflow_(fma2_fflags_lo_underflow_),
    .fma2_fflags_o_inexact_(fma2_fflags_lo_inexact_)
  );


  fpu_float_aux
  aux0
  (
    .fp_v_i(fp_v_i),
    .fpu_float_op_i(fpu_float_op_i),
    .fp_rs1_i(fp_rs1_i),
    .fp_rs2_i(fp_rs2_i),
    .fp_rm_i(fp_rm_i),
    .v_o(aux_v_lo),
    .result_o(aux_result_lo),
    .fflags_o_invalid_(aux_fflags_lo_invalid_),
    .fflags_o_div_zero_(aux_fflags_lo_div_zero_),
    .fflags_o_overflow_(aux_fflags_lo_overflow_),
    .fflags_o_underflow_(aux_fflags_lo_underflow_),
    .fflags_o_inexact_(aux_fflags_lo_inexact_)
  );

  assign N17 = (N0)? 1'b1 : 
               (N26)? 1'b1 : 
               (N16)? 1'b0 : 1'b0;
  assign N0 = N13;
  assign { N22, N21, N20, N19, N18 } = (N0)? fp_rd_i : 
                                       (N26)? imul_rd_i : 1'b0;
  assign N23 = (N1)? N17 : 
               (N2)? 1'b0 : 1'b0;
  assign N1 = N11;
  assign N2 = N12;
  assign N31 = (N3)? aux_v_lo : 
               (N4)? 1'b0 : 1'b0;
  assign N3 = N29;
  assign N4 = N30;
  assign N34 = (N5)? aux_v_r[0] : 
               (N6)? 1'b0 : 1'b0;
  assign N5 = N32;
  assign N6 = N33;
  assign { N36, N35 } = (N7)? { 1'b0, 1'b0 } : 
                        (N8)? { N34, N31 } : 1'b0;
  assign N7 = N28;
  assign N8 = N27;
  assign fp_result_o = (N9)? fma2_result_lo : 
                       (N10)? aux_result_r[65:33] : 1'b0;
  assign N9 = fma2_v_lo;
  assign N10 = N37;
  assign { fp_fflags_o_invalid_, fp_fflags_o_div_zero_, fp_fflags_o_overflow_, fp_fflags_o_underflow_, fp_fflags_o_inexact_ } = (N9)? { fma2_fflags_lo_invalid_, fma2_fflags_lo_div_zero_, fma2_fflags_lo_overflow_, fma2_fflags_lo_underflow_, fma2_fflags_lo_inexact_ } : 
                                                                                                                                (N10)? aux_fflags_r[9:5] : 1'b0;
  assign N11 = ~stall_fpu1_i;
  assign N12 = stall_fpu1_i;
  assign N13 = fp_v_i;
  assign N14 = imul_v_i;
  assign N15 = N14 | N13;
  assign N16 = ~N15;
  assign N24 = ~stall_fpu2_i;
  assign N25 = ~N13;
  assign N26 = N14 & N25;
  assign N27 = ~reset_i;
  assign N28 = reset_i;
  assign N29 = ~stall_fpu1_i;
  assign N30 = stall_fpu1_i;
  assign N32 = ~stall_fpu2_i;
  assign N33 = stall_fpu2_i;
  assign fpu1_v_r_o = fma1_v_lo | aux_v_r[0];
  assign fp_v_o = fma2_v_lo | aux_v_r[1];
  assign N37 = ~fma2_v_lo;

  always @(posedge clk_i) begin
    if(reset_i) begin
      fp_rd_o_4_sv2v_reg <= 1'b0;
      fp_rd_o_3_sv2v_reg <= 1'b0;
      fp_rd_o_2_sv2v_reg <= 1'b0;
      fp_rd_o_1_sv2v_reg <= 1'b0;
      fp_rd_o_0_sv2v_reg <= 1'b0;
    end else if(N24) begin
      fp_rd_o_4_sv2v_reg <= fpu1_rd_o[4];
      fp_rd_o_3_sv2v_reg <= fpu1_rd_o[3];
      fp_rd_o_2_sv2v_reg <= fpu1_rd_o[2];
      fp_rd_o_1_sv2v_reg <= fpu1_rd_o[1];
      fp_rd_o_0_sv2v_reg <= fpu1_rd_o[0];
    end 
    if(reset_i) begin
      fpu1_rd_o_4_sv2v_reg <= 1'b0;
      fpu1_rd_o_3_sv2v_reg <= 1'b0;
      fpu1_rd_o_2_sv2v_reg <= 1'b0;
      fpu1_rd_o_1_sv2v_reg <= 1'b0;
      fpu1_rd_o_0_sv2v_reg <= 1'b0;
    end else if(N23) begin
      fpu1_rd_o_4_sv2v_reg <= N22;
      fpu1_rd_o_3_sv2v_reg <= N21;
      fpu1_rd_o_2_sv2v_reg <= N20;
      fpu1_rd_o_1_sv2v_reg <= N19;
      fpu1_rd_o_0_sv2v_reg <= N18;
    end 
    if(N36) begin
      aux_fflags_r_9_sv2v_reg <= aux_fflags_r[4];
      aux_fflags_r_8_sv2v_reg <= aux_fflags_r[3];
      aux_fflags_r_7_sv2v_reg <= aux_fflags_r[2];
      aux_fflags_r_6_sv2v_reg <= aux_fflags_r[1];
      aux_fflags_r_5_sv2v_reg <= aux_fflags_r[0];
      aux_result_r_65_sv2v_reg <= aux_result_r[32];
      aux_result_r_64_sv2v_reg <= aux_result_r[31];
      aux_result_r_63_sv2v_reg <= aux_result_r[30];
      aux_result_r_62_sv2v_reg <= aux_result_r[29];
      aux_result_r_61_sv2v_reg <= aux_result_r[28];
      aux_result_r_60_sv2v_reg <= aux_result_r[27];
      aux_result_r_59_sv2v_reg <= aux_result_r[26];
      aux_result_r_58_sv2v_reg <= aux_result_r[25];
      aux_result_r_57_sv2v_reg <= aux_result_r[24];
      aux_result_r_56_sv2v_reg <= aux_result_r[23];
      aux_result_r_55_sv2v_reg <= aux_result_r[22];
      aux_result_r_54_sv2v_reg <= aux_result_r[21];
      aux_result_r_53_sv2v_reg <= aux_result_r[20];
      aux_result_r_52_sv2v_reg <= aux_result_r[19];
      aux_result_r_51_sv2v_reg <= aux_result_r[18];
      aux_result_r_50_sv2v_reg <= aux_result_r[17];
      aux_result_r_49_sv2v_reg <= aux_result_r[16];
      aux_result_r_48_sv2v_reg <= aux_result_r[15];
      aux_result_r_47_sv2v_reg <= aux_result_r[14];
      aux_result_r_46_sv2v_reg <= aux_result_r[13];
      aux_result_r_45_sv2v_reg <= aux_result_r[12];
      aux_result_r_44_sv2v_reg <= aux_result_r[11];
      aux_result_r_43_sv2v_reg <= aux_result_r[10];
      aux_result_r_42_sv2v_reg <= aux_result_r[9];
      aux_result_r_41_sv2v_reg <= aux_result_r[8];
      aux_result_r_40_sv2v_reg <= aux_result_r[7];
      aux_result_r_39_sv2v_reg <= aux_result_r[6];
      aux_result_r_38_sv2v_reg <= aux_result_r[5];
      aux_result_r_37_sv2v_reg <= aux_result_r[4];
      aux_result_r_36_sv2v_reg <= aux_result_r[3];
      aux_result_r_35_sv2v_reg <= aux_result_r[2];
      aux_result_r_34_sv2v_reg <= aux_result_r[1];
      aux_result_r_33_sv2v_reg <= aux_result_r[0];
    end 
    if(N35) begin
      aux_fflags_r_4_sv2v_reg <= aux_fflags_lo_invalid_;
      aux_fflags_r_3_sv2v_reg <= aux_fflags_lo_div_zero_;
      aux_fflags_r_2_sv2v_reg <= aux_fflags_lo_overflow_;
      aux_fflags_r_1_sv2v_reg <= aux_fflags_lo_underflow_;
      aux_fflags_r_0_sv2v_reg <= aux_fflags_lo_inexact_;
      aux_result_r_32_sv2v_reg <= aux_result_lo[32];
      aux_result_r_31_sv2v_reg <= aux_result_lo[31];
      aux_result_r_30_sv2v_reg <= aux_result_lo[30];
      aux_result_r_29_sv2v_reg <= aux_result_lo[29];
      aux_result_r_28_sv2v_reg <= aux_result_lo[28];
      aux_result_r_27_sv2v_reg <= aux_result_lo[27];
      aux_result_r_26_sv2v_reg <= aux_result_lo[26];
      aux_result_r_25_sv2v_reg <= aux_result_lo[25];
      aux_result_r_24_sv2v_reg <= aux_result_lo[24];
      aux_result_r_23_sv2v_reg <= aux_result_lo[23];
      aux_result_r_22_sv2v_reg <= aux_result_lo[22];
      aux_result_r_21_sv2v_reg <= aux_result_lo[21];
      aux_result_r_20_sv2v_reg <= aux_result_lo[20];
      aux_result_r_19_sv2v_reg <= aux_result_lo[19];
      aux_result_r_18_sv2v_reg <= aux_result_lo[18];
      aux_result_r_17_sv2v_reg <= aux_result_lo[17];
      aux_result_r_16_sv2v_reg <= aux_result_lo[16];
      aux_result_r_15_sv2v_reg <= aux_result_lo[15];
      aux_result_r_14_sv2v_reg <= aux_result_lo[14];
      aux_result_r_13_sv2v_reg <= aux_result_lo[13];
      aux_result_r_12_sv2v_reg <= aux_result_lo[12];
      aux_result_r_11_sv2v_reg <= aux_result_lo[11];
      aux_result_r_10_sv2v_reg <= aux_result_lo[10];
      aux_result_r_9_sv2v_reg <= aux_result_lo[9];
      aux_result_r_8_sv2v_reg <= aux_result_lo[8];
      aux_result_r_7_sv2v_reg <= aux_result_lo[7];
      aux_result_r_6_sv2v_reg <= aux_result_lo[6];
      aux_result_r_5_sv2v_reg <= aux_result_lo[5];
      aux_result_r_4_sv2v_reg <= aux_result_lo[4];
      aux_result_r_3_sv2v_reg <= aux_result_lo[3];
      aux_result_r_2_sv2v_reg <= aux_result_lo[2];
      aux_result_r_1_sv2v_reg <= aux_result_lo[1];
      aux_result_r_0_sv2v_reg <= aux_result_lo[0];
    end 
    if(reset_i) begin
      aux_v_r_1_sv2v_reg <= 1'b0;
    end else if(N32) begin
      aux_v_r_1_sv2v_reg <= aux_v_r[0];
    end 
    if(reset_i) begin
      aux_v_r_0_sv2v_reg <= 1'b0;
    end else if(N29) begin
      aux_v_r_0_sv2v_reg <= aux_v_lo;
    end 
  end


endmodule



module iNFromException_width32
(
  signedOut,
  isNaN,
  sign,
  out
);

  output [31:0] out;
  input signedOut;
  input isNaN;
  input sign;
  wire [31:0] out;
  wire out_30_,N0;
  assign out[0] = out_30_;
  assign out[1] = out_30_;
  assign out[2] = out_30_;
  assign out[3] = out_30_;
  assign out[4] = out_30_;
  assign out[5] = out_30_;
  assign out[6] = out_30_;
  assign out[7] = out_30_;
  assign out[8] = out_30_;
  assign out[9] = out_30_;
  assign out[10] = out_30_;
  assign out[11] = out_30_;
  assign out[12] = out_30_;
  assign out[13] = out_30_;
  assign out[14] = out_30_;
  assign out[15] = out_30_;
  assign out[16] = out_30_;
  assign out[17] = out_30_;
  assign out[18] = out_30_;
  assign out[19] = out_30_;
  assign out[20] = out_30_;
  assign out[21] = out_30_;
  assign out[22] = out_30_;
  assign out[23] = out_30_;
  assign out[24] = out_30_;
  assign out[25] = out_30_;
  assign out[26] = out_30_;
  assign out[27] = out_30_;
  assign out[28] = out_30_;
  assign out[29] = out_30_;
  assign out[30] = out_30_;
  assign out_30_ = isNaN | N0;
  assign N0 = ~sign;
  assign out[31] = signedOut ^ out_30_;

endmodule



module recFNToIN_expWidth8_sigWidth24_intWidth32
(
  control,
  in,
  roundingMode,
  signedOut,
  out,
  intExceptionFlags
);

  input [0:0] control;
  input [32:0] in;
  input [2:0] roundingMode;
  output [31:0] out;
  output [2:0] intExceptionFlags;
  input signedOut;
  wire [31:0] out,complUnroundedInt,roundedInt,excOut;
  wire [2:0] intExceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,isNaN,isInf,isZero,sign,magJustBelowOne,
  N12,N13,N14,N15,N16,N17,common_inexact,N18,roundIncr_near_even,
  roundIncr_near_maxMag,roundIncr,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,roundCarryBut2,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,common_overflow,N100,N101,N102,N103,N104,N105,
  N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255;
  wire [9:0] sExp;
  wire [24:0] sig;
  wire [54:0] shiftedSig;
  wire [0:0] alignedSig;

  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN
  (
    .in(in),
    .isNaN(isNaN),
    .isInf(isInf),
    .isZero(isZero),
    .sign(sign),
    .sExp(sExp),
    .sig(sig)
  );


  iNFromException_width32
  iNFromException
  (
    .signedOut(signedOut),
    .isNaN(isNaN),
    .sign(sign),
    .out(excOut)
  );

  assign N103 = ~sExp[4];
  assign N104 = ~sExp[3];
  assign N105 = ~sExp[2];
  assign N106 = ~sExp[1];
  assign N107 = ~sExp[0];
  assign N108 = sExp[6] | sExp[7];
  assign N109 = sExp[5] | N108;
  assign N110 = N103 | N109;
  assign N111 = N104 | N110;
  assign N112 = N105 | N111;
  assign N113 = N106 | N112;
  assign N114 = N107 | N113;
  assign N115 = ~N114;
  assign N116 = sExp[6] | sExp[7];
  assign N117 = sExp[5] | N116;
  assign N118 = N103 | N117;
  assign N119 = N104 | N118;
  assign N120 = N105 | N119;
  assign N121 = N106 | N120;
  assign N122 = sExp[0] | N121;
  assign N123 = ~N122;
  assign N124 = roundingMode[1] | roundingMode[2];
  assign N125 = roundingMode[0] | N124;
  assign N126 = ~N125;
  assign N127 = ~roundingMode[2];
  assign N128 = roundingMode[1] | N127;
  assign N129 = roundingMode[0] | N128;
  assign N130 = ~N129;
  assign N131 = ~roundingMode[1];
  assign N132 = N131 | roundingMode[2];
  assign N133 = roundingMode[0] | N132;
  assign N134 = ~N133;
  assign N135 = N131 | N127;
  assign N136 = roundingMode[0] | N135;
  assign N137 = ~N136;
  assign N138 = ~roundingMode[0];
  assign N139 = N138 | N132;
  assign N140 = ~N139;
  assign shiftedSig = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sExp[8:8], sig[22:0] } << { N16, N15, N14, N13, N12 };
  assign { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55 } = complUnroundedInt + 1'b1;
  assign { N16, N15, N14, N13, N12 } = (N0)? sExp[4:0] : 
                                       (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = sExp[8];
  assign N1 = N141;
  assign common_inexact = (N0)? N17 : 
                          (N1)? N18 : 1'b0;
  assign complUnroundedInt = (N2)? { N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52 } : 
                             (N3)? shiftedSig[54:23] : 1'b0;
  assign N2 = N20;
  assign N3 = N19;
  assign { roundedInt[31:1], N87 } = (N4)? { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55 } : 
                                     (N54)? complUnroundedInt : 1'b0;
  assign N4 = N53;
  assign N94 = (N5)? N92 : 
               (N6)? N93 : 1'b0;
  assign N5 = N91;
  assign N6 = N90;
  assign N96 = (N7)? N94 : 
               (N8)? N95 : 1'b0;
  assign N7 = N89;
  assign N8 = N88;
  assign N99 = (N9)? 1'b1 : 
               (N10)? N96 : 1'b0;
  assign N9 = N97;
  assign N10 = N98;
  assign common_overflow = (N0)? N99 : 
                           (N1)? N100 : 1'b0;
  assign out = (N11)? excOut : 
               (N102)? roundedInt : 1'b0;
  assign N11 = N101;
  assign magJustBelowOne = N141 & N148;
  assign N141 = ~sExp[8];
  assign N148 = N147 & sExp[0];
  assign N147 = N146 & sExp[1];
  assign N146 = N145 & sExp[2];
  assign N145 = N144 & sExp[3];
  assign N144 = N143 & sExp[4];
  assign N143 = N142 & sExp[5];
  assign N142 = sExp[7] & sExp[6];
  assign alignedSig[0] = N168 | shiftedSig[0];
  assign N168 = N167 | shiftedSig[1];
  assign N167 = N166 | shiftedSig[2];
  assign N166 = N165 | shiftedSig[3];
  assign N165 = N164 | shiftedSig[4];
  assign N164 = N163 | shiftedSig[5];
  assign N163 = N162 | shiftedSig[6];
  assign N162 = N161 | shiftedSig[7];
  assign N161 = N160 | shiftedSig[8];
  assign N160 = N159 | shiftedSig[9];
  assign N159 = N158 | shiftedSig[10];
  assign N158 = N157 | shiftedSig[11];
  assign N157 = N156 | shiftedSig[12];
  assign N156 = N155 | shiftedSig[13];
  assign N155 = N154 | shiftedSig[14];
  assign N154 = N153 | shiftedSig[15];
  assign N153 = N152 | shiftedSig[16];
  assign N152 = N151 | shiftedSig[17];
  assign N151 = N150 | shiftedSig[18];
  assign N150 = N149 | shiftedSig[19];
  assign N149 = shiftedSig[21] | shiftedSig[20];
  assign N17 = shiftedSig[22] | alignedSig[0];
  assign N18 = ~isZero;
  assign roundIncr_near_even = N172 | N174;
  assign N172 = sExp[8] & N171;
  assign N171 = N169 | N170;
  assign N169 = shiftedSig[23] & shiftedSig[22];
  assign N170 = shiftedSig[22] & alignedSig[0];
  assign N174 = magJustBelowOne & N173;
  assign N173 = shiftedSig[22] | alignedSig[0];
  assign roundIncr_near_maxMag = N175 | magJustBelowOne;
  assign N175 = sExp[8] & shiftedSig[22];
  assign roundIncr = N182 | N185;
  assign N182 = N178 | N181;
  assign N178 = N176 | N177;
  assign N176 = N126 & roundIncr_near_even;
  assign N177 = N130 & roundIncr_near_maxMag;
  assign N181 = N179 & N180;
  assign N179 = N134 | N137;
  assign N180 = sign & common_inexact;
  assign N185 = N140 & N184;
  assign N184 = N183 & common_inexact;
  assign N183 = ~sign;
  assign N19 = ~sign;
  assign N20 = sign;
  assign N21 = ~shiftedSig[54];
  assign N22 = ~shiftedSig[53];
  assign N23 = ~shiftedSig[52];
  assign N24 = ~shiftedSig[51];
  assign N25 = ~shiftedSig[50];
  assign N26 = ~shiftedSig[49];
  assign N27 = ~shiftedSig[48];
  assign N28 = ~shiftedSig[47];
  assign N29 = ~shiftedSig[46];
  assign N30 = ~shiftedSig[45];
  assign N31 = ~shiftedSig[44];
  assign N32 = ~shiftedSig[43];
  assign N33 = ~shiftedSig[42];
  assign N34 = ~shiftedSig[41];
  assign N35 = ~shiftedSig[40];
  assign N36 = ~shiftedSig[39];
  assign N37 = ~shiftedSig[38];
  assign N38 = ~shiftedSig[37];
  assign N39 = ~shiftedSig[36];
  assign N40 = ~shiftedSig[35];
  assign N41 = ~shiftedSig[34];
  assign N42 = ~shiftedSig[33];
  assign N43 = ~shiftedSig[32];
  assign N44 = ~shiftedSig[31];
  assign N45 = ~shiftedSig[30];
  assign N46 = ~shiftedSig[29];
  assign N47 = ~shiftedSig[28];
  assign N48 = ~shiftedSig[27];
  assign N49 = ~shiftedSig[26];
  assign N50 = ~shiftedSig[25];
  assign N51 = ~shiftedSig[24];
  assign N52 = ~shiftedSig[23];
  assign N53 = roundIncr ^ sign;
  assign N54 = ~N53;
  assign roundedInt[0] = N87 | N186;
  assign N186 = N137 & common_inexact;
  assign roundCarryBut2 = N215 & roundIncr;
  assign N215 = N214 & shiftedSig[23];
  assign N214 = N213 & shiftedSig[24];
  assign N213 = N212 & shiftedSig[25];
  assign N212 = N211 & shiftedSig[26];
  assign N211 = N210 & shiftedSig[27];
  assign N210 = N209 & shiftedSig[28];
  assign N209 = N208 & shiftedSig[29];
  assign N208 = N207 & shiftedSig[30];
  assign N207 = N206 & shiftedSig[31];
  assign N206 = N205 & shiftedSig[32];
  assign N205 = N204 & shiftedSig[33];
  assign N204 = N203 & shiftedSig[34];
  assign N203 = N202 & shiftedSig[35];
  assign N202 = N201 & shiftedSig[36];
  assign N201 = N200 & shiftedSig[37];
  assign N200 = N199 & shiftedSig[38];
  assign N199 = N198 & shiftedSig[39];
  assign N198 = N197 & shiftedSig[40];
  assign N197 = N196 & shiftedSig[41];
  assign N196 = N195 & shiftedSig[42];
  assign N195 = N194 & shiftedSig[43];
  assign N194 = N193 & shiftedSig[44];
  assign N193 = N192 & shiftedSig[45];
  assign N192 = N191 & shiftedSig[46];
  assign N191 = N190 & shiftedSig[47];
  assign N190 = N189 & shiftedSig[48];
  assign N189 = N188 & shiftedSig[49];
  assign N188 = N187 & shiftedSig[50];
  assign N187 = shiftedSig[52] & shiftedSig[51];
  assign N88 = ~signedOut;
  assign N89 = signedOut;
  assign N90 = ~sign;
  assign N91 = sign;
  assign N92 = N115 & N246;
  assign N246 = N245 | roundIncr;
  assign N245 = N244 | shiftedSig[23];
  assign N244 = N243 | shiftedSig[24];
  assign N243 = N242 | shiftedSig[25];
  assign N242 = N241 | shiftedSig[26];
  assign N241 = N240 | shiftedSig[27];
  assign N240 = N239 | shiftedSig[28];
  assign N239 = N238 | shiftedSig[29];
  assign N238 = N237 | shiftedSig[30];
  assign N237 = N236 | shiftedSig[31];
  assign N236 = N235 | shiftedSig[32];
  assign N235 = N234 | shiftedSig[33];
  assign N234 = N233 | shiftedSig[34];
  assign N233 = N232 | shiftedSig[35];
  assign N232 = N231 | shiftedSig[36];
  assign N231 = N230 | shiftedSig[37];
  assign N230 = N229 | shiftedSig[38];
  assign N229 = N228 | shiftedSig[39];
  assign N228 = N227 | shiftedSig[40];
  assign N227 = N226 | shiftedSig[41];
  assign N226 = N225 | shiftedSig[42];
  assign N225 = N224 | shiftedSig[43];
  assign N224 = N223 | shiftedSig[44];
  assign N223 = N222 | shiftedSig[45];
  assign N222 = N221 | shiftedSig[46];
  assign N221 = N220 | shiftedSig[47];
  assign N220 = N219 | shiftedSig[48];
  assign N219 = N218 | shiftedSig[49];
  assign N218 = N217 | shiftedSig[50];
  assign N217 = N216 | shiftedSig[51];
  assign N216 = shiftedSig[53] | shiftedSig[52];
  assign N93 = N115 | N247;
  assign N247 = N123 & roundCarryBut2;
  assign N95 = sign | N249;
  assign N249 = N248 & roundCarryBut2;
  assign N248 = N115 & shiftedSig[53];
  assign N97 = N250 | sExp[5];
  assign N250 = sExp[7] | sExp[6];
  assign N98 = ~N97;
  assign N100 = N252 & roundIncr;
  assign N252 = N251 & sign;
  assign N251 = ~signedOut;
  assign intExceptionFlags[2] = isNaN | isInf;
  assign intExceptionFlags[1] = N253 & common_overflow;
  assign N253 = ~intExceptionFlags[2];
  assign intExceptionFlags[0] = N255 & common_inexact;
  assign N255 = N253 & N254;
  assign N254 = ~common_overflow;
  assign N101 = intExceptionFlags[2] | common_overflow;
  assign N102 = ~N101;

endmodule



module fpu_int_fclass_exp_width_p8_sig_width_p24
(
  i,
  o
);

  input [32:0] i;
  output [9:0] o;
  wire [9:0] o,exp;
  wire is_nan,is_inf,is_zero,sign,N0,is_subnormal,is_normal,N1,N2,N3,N4,N5,N6,N7,N8,N9,
  N10,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,sv2v_dc_6,sv2v_dc_7,
  sv2v_dc_8,sv2v_dc_9,sv2v_dc_10,sv2v_dc_11,sv2v_dc_12,sv2v_dc_13,sv2v_dc_14,sv2v_dc_15,
  sv2v_dc_16,sv2v_dc_17,sv2v_dc_18,sv2v_dc_19,sv2v_dc_20,sv2v_dc_21,sv2v_dc_22,
  sv2v_dc_23,sv2v_dc_24,sv2v_dc_25;

  recFNToRawFN_expWidth8_sigWidth24
  raw0
  (
    .in(i),
    .isNaN(is_nan),
    .isInf(is_inf),
    .isZero(is_zero),
    .sign(sign),
    .sExp(exp),
    .sig({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6, sv2v_dc_7, sv2v_dc_8, sv2v_dc_9, sv2v_dc_10, sv2v_dc_11, sv2v_dc_12, sv2v_dc_13, sv2v_dc_14, sv2v_dc_15, sv2v_dc_16, sv2v_dc_17, sv2v_dc_18, sv2v_dc_19, sv2v_dc_20, sv2v_dc_21, sv2v_dc_22, sv2v_dc_23, sv2v_dc_24, sv2v_dc_25 })
  );

  assign N0 = exp < { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign is_subnormal = N4 & N5;
  assign N4 = N2 & N3;
  assign N2 = N0 & N1;
  assign N1 = ~is_nan;
  assign N3 = ~is_inf;
  assign N5 = ~is_zero;
  assign is_normal = ~N8;
  assign N8 = N7 | is_nan;
  assign N7 = N6 | is_zero;
  assign N6 = is_subnormal | is_inf;
  assign o[0] = sign & is_inf;
  assign o[1] = sign & is_normal;
  assign o[2] = sign & is_subnormal;
  assign o[3] = sign & is_zero;
  assign o[4] = N9 & is_zero;
  assign N9 = ~sign;
  assign o[5] = N9 & is_subnormal;
  assign o[6] = N9 & is_normal;
  assign o[7] = N9 & is_inf;
  assign o[8] = is_nan & N10;
  assign N10 = ~i[22];
  assign o[9] = is_nan & i[22];

endmodule



module fpu_int
(
  fp_rs1_i,
  fp_rs2_i,
  fpu_int_op_i,
  fp_rm_i,
  result_o,
  fflags_o_invalid_,
  fflags_o_div_zero_,
  fflags_o_overflow_,
  fflags_o_underflow_,
  fflags_o_inexact_
);

  input [32:0] fp_rs1_i;
  input [32:0] fp_rs2_i;
  input [2:0] fpu_int_op_i;
  input [2:0] fp_rm_i;
  output [31:0] result_o;
  output fflags_o_invalid_;
  output fflags_o_div_zero_;
  output fflags_o_overflow_;
  output fflags_o_underflow_;
  output fflags_o_inexact_;
  wire [31:0] result_o,f2i_result_lo,fp_rs1_fn;
  wire fflags_o_invalid_,fflags_o_div_zero_,fflags_o_overflow_,fflags_o_underflow_,
  fflags_o_inexact_,N0,N1,N2,cmp_signaling_li,cmp_lt_lo,cmp_eq_lo,cmp_unordered_lo,
  cmp_fflags_lo_invalid_,cmp_fflags_lo_div_zero_,cmp_fflags_lo_overflow_,
  cmp_fflags_lo_underflow_,cmp_fflags_lo_inexact_,cmp_result,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,f2i_fflags_lo_invalid_,f2i_fflags_lo_overflow_,f2i_fflags_lo_inexact_,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43;
  wire [9:0] fclass_result_lo;

  compareRecFN_expWidth8_sigWidth24
  cmp0
  (
    .a(fp_rs1_i),
    .b(fp_rs2_i),
    .signaling(cmp_signaling_li),
    .lt(cmp_lt_lo),
    .eq(cmp_eq_lo),
    .unordered(cmp_unordered_lo),
    .exceptionFlags({ cmp_fflags_lo_invalid_, cmp_fflags_lo_div_zero_, cmp_fflags_lo_overflow_, cmp_fflags_lo_underflow_, cmp_fflags_lo_inexact_ })
  );


  recFNToIN_expWidth8_sigWidth24_intWidth32
  f2i
  (
    .control(1'b1),
    .in(fp_rs1_i),
    .roundingMode(fp_rm_i),
    .signedOut(N33),
    .out(f2i_result_lo),
    .intExceptionFlags({ f2i_fflags_lo_invalid_, f2i_fflags_lo_overflow_, f2i_fflags_lo_inexact_ })
  );


  fpu_int_fclass_exp_width_p8_sig_width_p24
  fclass0
  (
    .i(fp_rs1_i),
    .o(fclass_result_lo)
  );


  recFNToFN_expWidth8_sigWidth24
  toFN0
  (
    .in(fp_rs1_i),
    .out(fp_rs1_fn)
  );

  assign N25 = ~fpu_int_op_i[2];
  assign N26 = ~fpu_int_op_i[0];
  assign N27 = fpu_int_op_i[1] | N25;
  assign N28 = N26 | N27;
  assign N29 = ~N28;
  assign N30 = ~fpu_int_op_i[1];
  assign N31 = N30 | fpu_int_op_i[2];
  assign N32 = N26 | N31;
  assign N33 = ~N32;
  assign N34 = fpu_int_op_i[0] | N27;
  assign N35 = ~N34;
  assign N36 = fpu_int_op_i[1] | fpu_int_op_i[2];
  assign N37 = N26 | N36;
  assign N38 = ~N37;
  assign N39 = fpu_int_op_i[0] | N36;
  assign N40 = ~N39;
  assign N41 = fpu_int_op_i[0] | N31;
  assign N42 = ~N41;
  assign cmp_result = (N0)? 1'b0 : 
                      (N9)? cmp_lt_lo : 
                      (N11)? N7 : 
                      (N13)? cmp_eq_lo : 
                      (N6)? 1'b0 : 1'b0;
  assign N0 = cmp_unordered_lo;
  assign result_o = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cmp_result } : 
                    (N21)? f2i_result_lo : 
                    (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fclass_result_lo } : 
                    (N18)? fp_rs1_fn : 1'b0;
  assign N1 = N14;
  assign { fflags_o_invalid_, fflags_o_overflow_, fflags_o_inexact_ } = (N1)? { cmp_fflags_lo_invalid_, cmp_fflags_lo_overflow_, cmp_fflags_lo_inexact_ } : 
                                                                        (N21)? { f2i_fflags_lo_invalid_, f2i_fflags_lo_overflow_, f2i_fflags_lo_inexact_ } : 
                                                                        (N19)? { 1'b0, 1'b0, 1'b0 } : 
                                                                        (N2)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = 1'b0;
  assign { fflags_o_div_zero_, fflags_o_underflow_ } = (N1)? { cmp_fflags_lo_div_zero_, cmp_fflags_lo_underflow_ } : 
                                                       (N20)? { 1'b0, 1'b0 } : 
                                                       (N2)? { 1'b0, 1'b0 } : 
                                                       (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign cmp_signaling_li = N42 | N38;
  assign N3 = N42 | cmp_unordered_lo;
  assign N4 = N38 | N3;
  assign N5 = N40 | N4;
  assign N6 = ~N5;
  assign N7 = cmp_lt_lo | cmp_eq_lo;
  assign N8 = ~cmp_unordered_lo;
  assign N9 = N42 & N8;
  assign N10 = N8 & N41;
  assign N11 = N38 & N10;
  assign N12 = N10 & N37;
  assign N13 = N40 & N12;
  assign N14 = N43 | N40;
  assign N43 = N42 | N38;
  assign N15 = N33 | N35;
  assign N16 = N15 | N14;
  assign N17 = N29 | N16;
  assign N18 = ~N17;
  assign N19 = ~N16;
  assign N20 = ~N14;
  assign N21 = N15 & N20;
  assign N22 = ~N15;
  assign N23 = N20 & N22;
  assign N24 = N29 & N23;

endmodule



module divSqrtRecFNToRaw_small_expWidth8_sigWidth24_options0
(
  nReset,
  clock,
  control,
  inReady,
  inValid,
  sqrtOp,
  a,
  b,
  roundingMode,
  outValid,
  sqrtOpOut,
  roundingModeOut,
  invalidExc,
  infiniteExc,
  out_isNaN,
  out_isInf,
  out_isZero,
  out_sign,
  out_sExp,
  out_sig
);

  input [0:0] control;
  input [32:0] a;
  input [32:0] b;
  input [2:0] roundingMode;
  output [2:0] roundingModeOut;
  output [9:0] out_sExp;
  output [26:0] out_sig;
  input nReset;
  input clock;
  input inValid;
  input sqrtOp;
  output inReady;
  output outValid;
  output sqrtOpOut;
  output invalidExc;
  output infiniteExc;
  output out_isNaN;
  output out_isInf;
  output out_isZero;
  output out_sign;
  wire [2:0] roundingModeOut;
  wire [9:0] out_sExp,sExpA_S,sExpB_S;
  wire [26:0] out_sig;
  wire inReady,outValid,sqrtOpOut,invalidExc,infiniteExc,out_isNaN,out_isInf,
  out_isZero,out_sign,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,isNaNA_S,
  isInfA_S,isZeroA_S,signA_S,isSigNaNA_S,isNaNB_S,isInfB_S,isZeroB_S,signB_S,
  isSigNaNB_S,notSigNaNIn_invalidExc_S_div,notSigNaNIn_invalidExc_S_sqrt,N17,N18,
  majorExc_S,N19,N20,isNaN_S,N21,isInf_S,N22,isZero_S,N23,sign_S,specialCaseA_S,
  specialCaseB_S,normalCase_S_div,normalCase_S_sqrt,normalCase_S,N24,N25,N26,N27,N28,N29,N30,
  N31,N32,N33,evenSqrt_S,oddSqrt_S,entering,entering_normalCase,skipCycle2,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,majorExc_Z,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,newBit,N268,
  N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,
  N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,
  N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,
  N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,sv2v_dc_1,sv2v_dc_2;
  wire [24:0] sigA_S,sigB_S,bitMask;
  wire [10:0] sExpQuot_S_div;
  wire [9:6] sSatExpQuot_S_div;
  wire [4:0] cycleNum;
  wire [22:0] fractB_Z;
  wire [1:0] decHiSigA_S;
  wire [25:0] rem_Z,trialTerm;
  wire [26:1] rem;
  wire [27:0] trialRem;
  reg cycleNum_4_sv2v_reg,cycleNum_3_sv2v_reg,cycleNum_2_sv2v_reg,cycleNum_1_sv2v_reg,
  cycleNum_0_sv2v_reg,fractB_Z_22_sv2v_reg,fractB_Z_21_sv2v_reg,
  fractB_Z_20_sv2v_reg,fractB_Z_19_sv2v_reg,fractB_Z_18_sv2v_reg,fractB_Z_17_sv2v_reg,
  fractB_Z_16_sv2v_reg,fractB_Z_15_sv2v_reg,fractB_Z_14_sv2v_reg,fractB_Z_13_sv2v_reg,
  fractB_Z_12_sv2v_reg,fractB_Z_11_sv2v_reg,fractB_Z_10_sv2v_reg,fractB_Z_9_sv2v_reg,
  fractB_Z_8_sv2v_reg,fractB_Z_7_sv2v_reg,fractB_Z_6_sv2v_reg,fractB_Z_5_sv2v_reg,
  fractB_Z_4_sv2v_reg,fractB_Z_3_sv2v_reg,fractB_Z_2_sv2v_reg,fractB_Z_1_sv2v_reg,
  fractB_Z_0_sv2v_reg,sqrtOpOut_sv2v_reg,majorExc_Z_sv2v_reg,out_isNaN_sv2v_reg,
  out_isInf_sv2v_reg,out_isZero_sv2v_reg,out_sign_sv2v_reg,out_sExp_9_sv2v_reg,
  out_sExp_8_sv2v_reg,out_sExp_7_sv2v_reg,out_sExp_6_sv2v_reg,out_sExp_5_sv2v_reg,
  out_sExp_4_sv2v_reg,out_sExp_3_sv2v_reg,out_sExp_2_sv2v_reg,out_sExp_1_sv2v_reg,
  out_sExp_0_sv2v_reg,roundingModeOut_2_sv2v_reg,roundingModeOut_1_sv2v_reg,
  roundingModeOut_0_sv2v_reg,out_sig_0_sv2v_reg,rem_Z_25_sv2v_reg,rem_Z_24_sv2v_reg,
  rem_Z_23_sv2v_reg,rem_Z_22_sv2v_reg,rem_Z_21_sv2v_reg,rem_Z_20_sv2v_reg,rem_Z_19_sv2v_reg,
  rem_Z_18_sv2v_reg,rem_Z_17_sv2v_reg,rem_Z_16_sv2v_reg,rem_Z_15_sv2v_reg,
  rem_Z_14_sv2v_reg,rem_Z_13_sv2v_reg,rem_Z_12_sv2v_reg,rem_Z_11_sv2v_reg,rem_Z_10_sv2v_reg,
  rem_Z_9_sv2v_reg,rem_Z_8_sv2v_reg,rem_Z_7_sv2v_reg,rem_Z_6_sv2v_reg,
  rem_Z_5_sv2v_reg,rem_Z_4_sv2v_reg,rem_Z_3_sv2v_reg,rem_Z_2_sv2v_reg,rem_Z_1_sv2v_reg,
  rem_Z_0_sv2v_reg,out_sig_26_sv2v_reg,out_sig_25_sv2v_reg,out_sig_24_sv2v_reg,
  out_sig_23_sv2v_reg,out_sig_22_sv2v_reg,out_sig_21_sv2v_reg,out_sig_20_sv2v_reg,
  out_sig_19_sv2v_reg,out_sig_18_sv2v_reg,out_sig_17_sv2v_reg,out_sig_16_sv2v_reg,
  out_sig_15_sv2v_reg,out_sig_14_sv2v_reg,out_sig_13_sv2v_reg,out_sig_12_sv2v_reg,
  out_sig_11_sv2v_reg,out_sig_10_sv2v_reg,out_sig_9_sv2v_reg,out_sig_8_sv2v_reg,
  out_sig_7_sv2v_reg,out_sig_6_sv2v_reg,out_sig_5_sv2v_reg,out_sig_4_sv2v_reg,out_sig_3_sv2v_reg,
  out_sig_2_sv2v_reg,out_sig_1_sv2v_reg;
  assign cycleNum[4] = cycleNum_4_sv2v_reg;
  assign cycleNum[3] = cycleNum_3_sv2v_reg;
  assign cycleNum[2] = cycleNum_2_sv2v_reg;
  assign cycleNum[1] = cycleNum_1_sv2v_reg;
  assign cycleNum[0] = cycleNum_0_sv2v_reg;
  assign fractB_Z[22] = fractB_Z_22_sv2v_reg;
  assign fractB_Z[21] = fractB_Z_21_sv2v_reg;
  assign fractB_Z[20] = fractB_Z_20_sv2v_reg;
  assign fractB_Z[19] = fractB_Z_19_sv2v_reg;
  assign fractB_Z[18] = fractB_Z_18_sv2v_reg;
  assign fractB_Z[17] = fractB_Z_17_sv2v_reg;
  assign fractB_Z[16] = fractB_Z_16_sv2v_reg;
  assign fractB_Z[15] = fractB_Z_15_sv2v_reg;
  assign fractB_Z[14] = fractB_Z_14_sv2v_reg;
  assign fractB_Z[13] = fractB_Z_13_sv2v_reg;
  assign fractB_Z[12] = fractB_Z_12_sv2v_reg;
  assign fractB_Z[11] = fractB_Z_11_sv2v_reg;
  assign fractB_Z[10] = fractB_Z_10_sv2v_reg;
  assign fractB_Z[9] = fractB_Z_9_sv2v_reg;
  assign fractB_Z[8] = fractB_Z_8_sv2v_reg;
  assign fractB_Z[7] = fractB_Z_7_sv2v_reg;
  assign fractB_Z[6] = fractB_Z_6_sv2v_reg;
  assign fractB_Z[5] = fractB_Z_5_sv2v_reg;
  assign fractB_Z[4] = fractB_Z_4_sv2v_reg;
  assign fractB_Z[3] = fractB_Z_3_sv2v_reg;
  assign fractB_Z[2] = fractB_Z_2_sv2v_reg;
  assign fractB_Z[1] = fractB_Z_1_sv2v_reg;
  assign fractB_Z[0] = fractB_Z_0_sv2v_reg;
  assign sqrtOpOut = sqrtOpOut_sv2v_reg;
  assign majorExc_Z = majorExc_Z_sv2v_reg;
  assign out_isNaN = out_isNaN_sv2v_reg;
  assign out_isInf = out_isInf_sv2v_reg;
  assign out_isZero = out_isZero_sv2v_reg;
  assign out_sign = out_sign_sv2v_reg;
  assign out_sExp[9] = out_sExp_9_sv2v_reg;
  assign out_sExp[8] = out_sExp_8_sv2v_reg;
  assign out_sExp[7] = out_sExp_7_sv2v_reg;
  assign out_sExp[6] = out_sExp_6_sv2v_reg;
  assign out_sExp[5] = out_sExp_5_sv2v_reg;
  assign out_sExp[4] = out_sExp_4_sv2v_reg;
  assign out_sExp[3] = out_sExp_3_sv2v_reg;
  assign out_sExp[2] = out_sExp_2_sv2v_reg;
  assign out_sExp[1] = out_sExp_1_sv2v_reg;
  assign out_sExp[0] = out_sExp_0_sv2v_reg;
  assign roundingModeOut[2] = roundingModeOut_2_sv2v_reg;
  assign roundingModeOut[1] = roundingModeOut_1_sv2v_reg;
  assign roundingModeOut[0] = roundingModeOut_0_sv2v_reg;
  assign out_sig[0] = out_sig_0_sv2v_reg;
  assign rem_Z[25] = rem_Z_25_sv2v_reg;
  assign rem_Z[24] = rem_Z_24_sv2v_reg;
  assign rem_Z[23] = rem_Z_23_sv2v_reg;
  assign rem_Z[22] = rem_Z_22_sv2v_reg;
  assign rem_Z[21] = rem_Z_21_sv2v_reg;
  assign rem_Z[20] = rem_Z_20_sv2v_reg;
  assign rem_Z[19] = rem_Z_19_sv2v_reg;
  assign rem_Z[18] = rem_Z_18_sv2v_reg;
  assign rem_Z[17] = rem_Z_17_sv2v_reg;
  assign rem_Z[16] = rem_Z_16_sv2v_reg;
  assign rem_Z[15] = rem_Z_15_sv2v_reg;
  assign rem_Z[14] = rem_Z_14_sv2v_reg;
  assign rem_Z[13] = rem_Z_13_sv2v_reg;
  assign rem_Z[12] = rem_Z_12_sv2v_reg;
  assign rem_Z[11] = rem_Z_11_sv2v_reg;
  assign rem_Z[10] = rem_Z_10_sv2v_reg;
  assign rem_Z[9] = rem_Z_9_sv2v_reg;
  assign rem_Z[8] = rem_Z_8_sv2v_reg;
  assign rem_Z[7] = rem_Z_7_sv2v_reg;
  assign rem_Z[6] = rem_Z_6_sv2v_reg;
  assign rem_Z[5] = rem_Z_5_sv2v_reg;
  assign rem_Z[4] = rem_Z_4_sv2v_reg;
  assign rem_Z[3] = rem_Z_3_sv2v_reg;
  assign rem_Z[2] = rem_Z_2_sv2v_reg;
  assign rem_Z[1] = rem_Z_1_sv2v_reg;
  assign rem_Z[0] = rem_Z_0_sv2v_reg;
  assign out_sig[26] = out_sig_26_sv2v_reg;
  assign out_sig[25] = out_sig_25_sv2v_reg;
  assign out_sig[24] = out_sig_24_sv2v_reg;
  assign out_sig[23] = out_sig_23_sv2v_reg;
  assign out_sig[22] = out_sig_22_sv2v_reg;
  assign out_sig[21] = out_sig_21_sv2v_reg;
  assign out_sig[20] = out_sig_20_sv2v_reg;
  assign out_sig[19] = out_sig_19_sv2v_reg;
  assign out_sig[18] = out_sig_18_sv2v_reg;
  assign out_sig[17] = out_sig_17_sv2v_reg;
  assign out_sig[16] = out_sig_16_sv2v_reg;
  assign out_sig[15] = out_sig_15_sv2v_reg;
  assign out_sig[14] = out_sig_14_sv2v_reg;
  assign out_sig[13] = out_sig_13_sv2v_reg;
  assign out_sig[12] = out_sig_12_sv2v_reg;
  assign out_sig[11] = out_sig_11_sv2v_reg;
  assign out_sig[10] = out_sig_10_sv2v_reg;
  assign out_sig[9] = out_sig_9_sv2v_reg;
  assign out_sig[8] = out_sig_8_sv2v_reg;
  assign out_sig[7] = out_sig_7_sv2v_reg;
  assign out_sig[6] = out_sig_6_sv2v_reg;
  assign out_sig[5] = out_sig_5_sv2v_reg;
  assign out_sig[4] = out_sig_4_sv2v_reg;
  assign out_sig[3] = out_sig_3_sv2v_reg;
  assign out_sig[2] = out_sig_2_sv2v_reg;
  assign out_sig[1] = out_sig_1_sv2v_reg;

  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN_a
  (
    .in(a),
    .isNaN(isNaNA_S),
    .isInf(isInfA_S),
    .isZero(isZeroA_S),
    .sign(signA_S),
    .sExp(sExpA_S),
    .sig(sigA_S)
  );


  isSigNaNRecFN_expWidth8_sigWidth24
  isSigNaN_a
  (
    .in(a),
    .isSigNaN(isSigNaNA_S)
  );


  recFNToRawFN_expWidth8_sigWidth24
  recFNToRawFN_b
  (
    .in(b),
    .isNaN(isNaNB_S),
    .isInf(isInfB_S),
    .isZero(isZeroB_S),
    .sign(signB_S),
    .sExp(sExpB_S),
    .sig(sigB_S)
  );


  isSigNaNRecFN_expWidth8_sigWidth24
  isSigNaN_b
  (
    .in(b),
    .isSigNaN(isSigNaNB_S)
  );

  assign N32 = $signed({ 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) <= $signed(sExpQuot_S_div);
  assign inReady = cycleNum <= 1'b1;
  assign { bitMask, sv2v_dc_1, sv2v_dc_2 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << cycleNum;
  assign newBit = $signed(1'b0) <= $signed(trialRem);
  assign N268 = cycleNum > { 1'b1, 1'b0 };
  assign N298 = $signed(trialRem) != $signed(1'b0);
  assign N360 = ~cycleNum[0];
  assign N361 = cycleNum[3] | cycleNum[4];
  assign N362 = cycleNum[2] | N361;
  assign N363 = cycleNum[1] | N362;
  assign N364 = N360 | N363;
  assign outValid = ~N364;
  assign N366 = cycleNum[3] | cycleNum[4];
  assign N367 = cycleNum[2] | N366;
  assign N368 = cycleNum[1] | N367;
  assign N369 = cycleNum[0] | N368;
  assign N370 = ~cycleNum[1];
  assign N371 = cycleNum[3] | cycleNum[4];
  assign N372 = cycleNum[2] | N371;
  assign N373 = N370 | N372;
  assign N374 = N360 | N373;
  assign N375 = ~N374;
  assign sExpQuot_S_div = sExpA_S + { sExpB_S[8:8], sExpB_S[8:8], sExpB_S[8:8], N24, N25, N26, N27, N28, N29, N30, N31 };
  assign decHiSigA_S = sigA_S[23:22] - 1'b1;
  assign { N71, N70, N69, N68, N67, N66, N65, N64, N63, N62 } = $signed(sExpA_S[9:1]) + $signed({ 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 });
  assign trialRem = { rem, 1'b0 } - trialTerm;
  assign { N48, N47, N46, N45, N44 } = cycleNum - 1'b1;
  assign majorExc_S = (N0)? N18 : 
                      (N1)? N19 : 1'b0;
  assign N0 = sqrtOp;
  assign N1 = N17;
  assign isNaN_S = (N0)? N20 : 
                   (N1)? N21 : 1'b0;
  assign isInf_S = (N0)? isInfA_S : 
                   (N1)? N22 : 1'b0;
  assign isZero_S = (N0)? isZeroA_S : 
                    (N1)? N23 : 1'b0;
  assign normalCase_S = (N0)? normalCase_S_sqrt : 
                        (N1)? normalCase_S_div : 1'b0;
  assign sSatExpQuot_S_div = (N2)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                             (N33)? sExpQuot_S_div[9:6] : 1'b0;
  assign N2 = N32;
  assign N38 = ~sExpA_S[0];
  assign N39 = (N0)? N38 : 
               (N1)? 1'b0 : 1'b0;
  assign { N41, N40 } = (N3)? { N17, N39 } : 
                        (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign N3 = entering_normalCase;
  assign N4 = N37;
  assign { N53, N52, N51, N50, N49 } = (N5)? { N48, N47, N46, N45, N44 } : 
                                       (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N42;
  assign { N81, N80, N79, N78, N77, N76, N75, N74, N73, N72 } = (N0)? { N71, N70, N69, N68, N67, N66, N65, N64, N63, N62 } : 
                                                                (N1)? { sSatExpQuot_S_div, sExpQuot_S_div[5:0] } : 1'b0;
  assign { N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85 } = (N6)? sigA_S : 
                                                                                                                                                     (N84)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N83;
  assign { N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112 } = (N7)? { decHiSigA_S, sigA_S[21:0] } : 
                                                                                                                                                              (N111)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N7 = N110;
  assign { N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137 } = (N8)? rem_Z : 
                                                                                                                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N136;
  assign N9 = inReady;
  assign { N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165 } = (N10)? sigB_S : 
                                                                                                                                                                    (N164)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = N163;
  assign { N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194 } = (N11)? fractB_Z : 
                                                                                                                                                        (N193)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N192;
  assign { N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, trialTerm[0:0] } = (N12)? { out_sig[25:25], N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, bitMask[0:0] } : 
                                                                                                                                                                                    (N218)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = N217;
  assign { N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271 } = (N13)? trialRem[25:0] : 
                                                                                                                                                                          (N14)? { rem[25:1], 1'b0 } : 1'b0;
  assign N13 = newBit;
  assign N14 = N270;
  assign N301 = (N15)? newBit : 
                (N300)? 1'b0 : 1'b0;
  assign N15 = N299;
  assign N305 = (N16)? newBit : 
                (N304)? 1'b0 : 1'b0;
  assign N16 = N303;
  assign { N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331 } = (N8)? { out_sig[26:26], N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330 } : 
                                                                                                                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign notSigNaNIn_invalidExc_S_div = N376 | N377;
  assign N376 = isZeroA_S & isZeroB_S;
  assign N377 = isInfA_S & isInfB_S;
  assign notSigNaNIn_invalidExc_S_sqrt = N380 & signA_S;
  assign N380 = N378 & N379;
  assign N378 = ~isNaNA_S;
  assign N379 = ~isZeroA_S;
  assign N17 = ~sqrtOp;
  assign N18 = isSigNaNA_S | notSigNaNIn_invalidExc_S_sqrt;
  assign N19 = N382 | N385;
  assign N382 = N381 | notSigNaNIn_invalidExc_S_div;
  assign N381 = isSigNaNA_S | isSigNaNB_S;
  assign N385 = N384 & isZeroB_S;
  assign N384 = N378 & N383;
  assign N383 = ~isInfA_S;
  assign N20 = isNaNA_S | notSigNaNIn_invalidExc_S_sqrt;
  assign N21 = N386 | notSigNaNIn_invalidExc_S_div;
  assign N386 = isNaNA_S | isNaNB_S;
  assign N22 = isInfA_S | isZeroB_S;
  assign N23 = isZeroA_S | isInfB_S;
  assign sign_S = signA_S ^ N387;
  assign N387 = N17 & signB_S;
  assign specialCaseA_S = N388 | isZeroA_S;
  assign N388 = isNaNA_S | isInfA_S;
  assign specialCaseB_S = N389 | isZeroB_S;
  assign N389 = isNaNB_S | isInfB_S;
  assign normalCase_S_div = N390 & N391;
  assign N390 = ~specialCaseA_S;
  assign N391 = ~specialCaseB_S;
  assign normalCase_S_sqrt = N390 & N392;
  assign N392 = ~signA_S;
  assign N24 = ~sExpB_S[7];
  assign N25 = ~sExpB_S[6];
  assign N26 = ~sExpB_S[5];
  assign N27 = ~sExpB_S[4];
  assign N28 = ~sExpB_S[3];
  assign N29 = ~sExpB_S[2];
  assign N30 = ~sExpB_S[1];
  assign N31 = ~sExpB_S[0];
  assign N33 = ~N32;
  assign evenSqrt_S = sqrtOp & N393;
  assign N393 = ~sExpA_S[0];
  assign oddSqrt_S = sqrtOp & sExpA_S[0];
  assign entering = inReady & inValid;
  assign entering_normalCase = entering & normalCase_S;
  assign skipCycle2 = N375 & out_sig[26];
  assign N34 = N369 | inValid;
  assign N35 = N60 & N34;
  assign N36 = entering & N394;
  assign N394 = ~normalCase_S;
  assign N37 = ~entering_normalCase;
  assign N42 = N369 & N395;
  assign N395 = ~skipCycle2;
  assign N43 = ~N42;
  assign N54 = N369 & skipCycle2;
  assign N55 = entering_normalCase | N53;
  assign N56 = entering_normalCase | N52;
  assign N57 = N41 | N50;
  assign N58 = N397 | N54;
  assign N397 = N396 | N49;
  assign N396 = N36 | N40;
  assign N59 = ~nReset;
  assign N60 = nReset;
  assign N61 = N60 & entering_normalCase;
  assign N82 = entering_normalCase & N17;
  assign N83 = inReady & N398;
  assign N398 = ~oddSqrt_S;
  assign N84 = ~N83;
  assign N110 = inReady & oddSqrt_S;
  assign N111 = ~N110;
  assign N136 = ~inReady;
  assign rem[26] = N135 | N162;
  assign rem[25] = N399 | N161;
  assign N399 = N109 | N134;
  assign rem[24] = N400 | N160;
  assign N400 = N108 | N133;
  assign rem[23] = N401 | N159;
  assign N401 = N107 | N132;
  assign rem[22] = N402 | N158;
  assign N402 = N106 | N131;
  assign rem[21] = N403 | N157;
  assign N403 = N105 | N130;
  assign rem[20] = N404 | N156;
  assign N404 = N104 | N129;
  assign rem[19] = N405 | N155;
  assign N405 = N103 | N128;
  assign rem[18] = N406 | N154;
  assign N406 = N102 | N127;
  assign rem[17] = N407 | N153;
  assign N407 = N101 | N126;
  assign rem[16] = N408 | N152;
  assign N408 = N100 | N125;
  assign rem[15] = N409 | N151;
  assign N409 = N99 | N124;
  assign rem[14] = N410 | N150;
  assign N410 = N98 | N123;
  assign rem[13] = N411 | N149;
  assign N411 = N97 | N122;
  assign rem[12] = N412 | N148;
  assign N412 = N96 | N121;
  assign rem[11] = N413 | N147;
  assign N413 = N95 | N120;
  assign rem[10] = N414 | N146;
  assign N414 = N94 | N119;
  assign rem[9] = N415 | N145;
  assign N415 = N93 | N118;
  assign rem[8] = N416 | N144;
  assign N416 = N92 | N117;
  assign rem[7] = N417 | N143;
  assign N417 = N91 | N116;
  assign rem[6] = N418 | N142;
  assign N418 = N90 | N115;
  assign rem[5] = N419 | N141;
  assign N419 = N89 | N114;
  assign rem[4] = N420 | N140;
  assign N420 = N88 | N113;
  assign rem[3] = N421 | N139;
  assign N421 = N87 | N112;
  assign rem[2] = N86 | N138;
  assign rem[1] = N85 | N137;
  assign N163 = inReady & N17;
  assign N164 = ~N163;
  assign N190 = inReady & evenSqrt_S;
  assign N191 = inReady & oddSqrt_S;
  assign N192 = N136 & N422;
  assign N422 = ~sqrtOpOut;
  assign N193 = ~N192;
  assign N217 = N136 & sqrtOpOut;
  assign N218 = ~N217;
  assign N219 = out_sig[24] | bitMask[24];
  assign N220 = out_sig[23] | bitMask[23];
  assign N221 = out_sig[22] | bitMask[22];
  assign N222 = out_sig[21] | bitMask[21];
  assign N223 = out_sig[20] | bitMask[20];
  assign N224 = out_sig[19] | bitMask[19];
  assign N225 = out_sig[18] | bitMask[18];
  assign N226 = out_sig[17] | bitMask[17];
  assign N227 = out_sig[16] | bitMask[16];
  assign N228 = out_sig[15] | bitMask[15];
  assign N229 = out_sig[14] | bitMask[14];
  assign N230 = out_sig[13] | bitMask[13];
  assign N231 = out_sig[12] | bitMask[12];
  assign N232 = out_sig[11] | bitMask[11];
  assign N233 = out_sig[10] | bitMask[10];
  assign N234 = out_sig[9] | bitMask[9];
  assign N235 = out_sig[8] | bitMask[8];
  assign N236 = out_sig[7] | bitMask[7];
  assign N237 = out_sig[6] | bitMask[6];
  assign N238 = out_sig[5] | bitMask[5];
  assign N239 = out_sig[4] | bitMask[4];
  assign N240 = out_sig[3] | bitMask[3];
  assign N241 = out_sig[2] | bitMask[2];
  assign N242 = out_sig[1] | bitMask[1];
  assign trialTerm[25] = N423 | N267;
  assign N423 = N189 | N191;
  assign trialTerm[24] = N425 | N266;
  assign N425 = N424 | N192;
  assign N424 = N188 | N190;
  assign trialTerm[23] = N427 | N265;
  assign N427 = N426 | N216;
  assign N426 = N187 | N191;
  assign trialTerm[22] = N428 | N264;
  assign N428 = N186 | N215;
  assign trialTerm[21] = N429 | N263;
  assign N429 = N185 | N214;
  assign trialTerm[20] = N430 | N262;
  assign N430 = N184 | N213;
  assign trialTerm[19] = N431 | N261;
  assign N431 = N183 | N212;
  assign trialTerm[18] = N432 | N260;
  assign N432 = N182 | N211;
  assign trialTerm[17] = N433 | N259;
  assign N433 = N181 | N210;
  assign trialTerm[16] = N434 | N258;
  assign N434 = N180 | N209;
  assign trialTerm[15] = N435 | N257;
  assign N435 = N179 | N208;
  assign trialTerm[14] = N436 | N256;
  assign N436 = N178 | N207;
  assign trialTerm[13] = N437 | N255;
  assign N437 = N177 | N206;
  assign trialTerm[12] = N438 | N254;
  assign N438 = N176 | N205;
  assign trialTerm[11] = N439 | N253;
  assign N439 = N175 | N204;
  assign trialTerm[10] = N440 | N252;
  assign N440 = N174 | N203;
  assign trialTerm[9] = N441 | N251;
  assign N441 = N173 | N202;
  assign trialTerm[8] = N442 | N250;
  assign N442 = N172 | N201;
  assign trialTerm[7] = N443 | N249;
  assign N443 = N171 | N200;
  assign trialTerm[6] = N444 | N248;
  assign N444 = N170 | N199;
  assign trialTerm[5] = N445 | N247;
  assign N445 = N169 | N198;
  assign trialTerm[4] = N446 | N246;
  assign N446 = N168 | N197;
  assign trialTerm[3] = N447 | N245;
  assign N447 = N167 | N196;
  assign trialTerm[2] = N448 | N244;
  assign N448 = N166 | N195;
  assign trialTerm[1] = N449 | N243;
  assign N449 = N165 | N194;
  assign N269 = entering_normalCase | N268;
  assign N270 = ~newBit;
  assign N297 = entering_normalCase | N450;
  assign N450 = N136 & newBit;
  assign N299 = inReady & N17;
  assign N300 = ~N299;
  assign N302 = inReady & sqrtOp;
  assign N303 = inReady & oddSqrt_S;
  assign N304 = ~N303;
  assign N306 = out_sig[25] | bitMask[24];
  assign N307 = out_sig[24] | bitMask[23];
  assign N308 = out_sig[23] | bitMask[22];
  assign N309 = out_sig[22] | bitMask[21];
  assign N310 = out_sig[21] | bitMask[20];
  assign N311 = out_sig[20] | bitMask[19];
  assign N312 = out_sig[19] | bitMask[18];
  assign N313 = out_sig[18] | bitMask[17];
  assign N314 = out_sig[17] | bitMask[16];
  assign N315 = out_sig[16] | bitMask[15];
  assign N316 = out_sig[15] | bitMask[14];
  assign N317 = out_sig[14] | bitMask[13];
  assign N318 = out_sig[13] | bitMask[12];
  assign N319 = out_sig[12] | bitMask[11];
  assign N320 = out_sig[11] | bitMask[10];
  assign N321 = out_sig[10] | bitMask[9];
  assign N322 = out_sig[9] | bitMask[8];
  assign N323 = out_sig[8] | bitMask[7];
  assign N324 = out_sig[7] | bitMask[6];
  assign N325 = out_sig[6] | bitMask[5];
  assign N326 = out_sig[5] | bitMask[4];
  assign N327 = out_sig[4] | bitMask[3];
  assign N328 = out_sig[3] | bitMask[2];
  assign N329 = out_sig[2] | bitMask[1];
  assign N330 = out_sig[1] | bitMask[0];
  assign N357 = N301 | N356;
  assign N358 = N302 | N355;
  assign N359 = N305 | N354;
  assign invalidExc = majorExc_Z & out_isNaN;
  assign infiniteExc = majorExc_Z & N451;
  assign N451 = ~out_isNaN;

  always @(posedge clock or posedge N59) begin
    if(N59) begin
      cycleNum_4_sv2v_reg <= 1'b0;
      cycleNum_3_sv2v_reg <= 1'b0;
      cycleNum_2_sv2v_reg <= 1'b0;
      cycleNum_1_sv2v_reg <= 1'b0;
      cycleNum_0_sv2v_reg <= 1'b0;
    end else if(N34) begin
      cycleNum_4_sv2v_reg <= N55;
      cycleNum_3_sv2v_reg <= N56;
      cycleNum_2_sv2v_reg <= N51;
      cycleNum_1_sv2v_reg <= N57;
      cycleNum_0_sv2v_reg <= N58;
    end 
  end


  always @(posedge clock) begin
    if(N59) begin
      fractB_Z_22_sv2v_reg <= 1'b0;
      fractB_Z_21_sv2v_reg <= 1'b0;
      fractB_Z_20_sv2v_reg <= 1'b0;
      fractB_Z_19_sv2v_reg <= 1'b0;
      fractB_Z_18_sv2v_reg <= 1'b0;
      fractB_Z_17_sv2v_reg <= 1'b0;
      fractB_Z_16_sv2v_reg <= 1'b0;
      fractB_Z_15_sv2v_reg <= 1'b0;
      fractB_Z_14_sv2v_reg <= 1'b0;
      fractB_Z_13_sv2v_reg <= 1'b0;
      fractB_Z_12_sv2v_reg <= 1'b0;
      fractB_Z_11_sv2v_reg <= 1'b0;
      fractB_Z_10_sv2v_reg <= 1'b0;
      fractB_Z_9_sv2v_reg <= 1'b0;
      fractB_Z_8_sv2v_reg <= 1'b0;
      fractB_Z_7_sv2v_reg <= 1'b0;
      fractB_Z_6_sv2v_reg <= 1'b0;
      fractB_Z_5_sv2v_reg <= 1'b0;
      fractB_Z_4_sv2v_reg <= 1'b0;
      fractB_Z_3_sv2v_reg <= 1'b0;
      fractB_Z_2_sv2v_reg <= 1'b0;
      fractB_Z_1_sv2v_reg <= 1'b0;
      fractB_Z_0_sv2v_reg <= 1'b0;
    end else if(N82) begin
      fractB_Z_22_sv2v_reg <= sigB_S[22];
      fractB_Z_21_sv2v_reg <= sigB_S[21];
      fractB_Z_20_sv2v_reg <= sigB_S[20];
      fractB_Z_19_sv2v_reg <= sigB_S[19];
      fractB_Z_18_sv2v_reg <= sigB_S[18];
      fractB_Z_17_sv2v_reg <= sigB_S[17];
      fractB_Z_16_sv2v_reg <= sigB_S[16];
      fractB_Z_15_sv2v_reg <= sigB_S[15];
      fractB_Z_14_sv2v_reg <= sigB_S[14];
      fractB_Z_13_sv2v_reg <= sigB_S[13];
      fractB_Z_12_sv2v_reg <= sigB_S[12];
      fractB_Z_11_sv2v_reg <= sigB_S[11];
      fractB_Z_10_sv2v_reg <= sigB_S[10];
      fractB_Z_9_sv2v_reg <= sigB_S[9];
      fractB_Z_8_sv2v_reg <= sigB_S[8];
      fractB_Z_7_sv2v_reg <= sigB_S[7];
      fractB_Z_6_sv2v_reg <= sigB_S[6];
      fractB_Z_5_sv2v_reg <= sigB_S[5];
      fractB_Z_4_sv2v_reg <= sigB_S[4];
      fractB_Z_3_sv2v_reg <= sigB_S[3];
      fractB_Z_2_sv2v_reg <= sigB_S[2];
      fractB_Z_1_sv2v_reg <= sigB_S[1];
      fractB_Z_0_sv2v_reg <= sigB_S[0];
    end 
    if(N59) begin
      sqrtOpOut_sv2v_reg <= 1'b0;
      majorExc_Z_sv2v_reg <= 1'b0;
      out_isNaN_sv2v_reg <= 1'b0;
      out_isInf_sv2v_reg <= 1'b0;
      out_isZero_sv2v_reg <= 1'b0;
      out_sign_sv2v_reg <= 1'b0;
    end else if(entering) begin
      sqrtOpOut_sv2v_reg <= sqrtOp;
      majorExc_Z_sv2v_reg <= majorExc_S;
      out_isNaN_sv2v_reg <= isNaN_S;
      out_isInf_sv2v_reg <= isInf_S;
      out_isZero_sv2v_reg <= isZero_S;
      out_sign_sv2v_reg <= sign_S;
    end 
    if(N59) begin
      out_sExp_9_sv2v_reg <= 1'b0;
      out_sExp_8_sv2v_reg <= 1'b0;
      out_sExp_7_sv2v_reg <= 1'b0;
      out_sExp_6_sv2v_reg <= 1'b0;
      out_sExp_5_sv2v_reg <= 1'b0;
      out_sExp_4_sv2v_reg <= 1'b0;
      out_sExp_3_sv2v_reg <= 1'b0;
      out_sExp_2_sv2v_reg <= 1'b0;
      out_sExp_1_sv2v_reg <= 1'b0;
      out_sExp_0_sv2v_reg <= 1'b0;
      roundingModeOut_2_sv2v_reg <= 1'b0;
      roundingModeOut_1_sv2v_reg <= 1'b0;
      roundingModeOut_0_sv2v_reg <= 1'b0;
    end else if(entering_normalCase) begin
      out_sExp_9_sv2v_reg <= N81;
      out_sExp_8_sv2v_reg <= N80;
      out_sExp_7_sv2v_reg <= N79;
      out_sExp_6_sv2v_reg <= N78;
      out_sExp_5_sv2v_reg <= N77;
      out_sExp_4_sv2v_reg <= N76;
      out_sExp_3_sv2v_reg <= N75;
      out_sExp_2_sv2v_reg <= N74;
      out_sExp_1_sv2v_reg <= N73;
      out_sExp_0_sv2v_reg <= N72;
      roundingModeOut_2_sv2v_reg <= roundingMode[2];
      roundingModeOut_1_sv2v_reg <= roundingMode[1];
      roundingModeOut_0_sv2v_reg <= roundingMode[0];
    end 
    if(N59) begin
      out_sig_0_sv2v_reg <= 1'b0;
      out_sig_26_sv2v_reg <= 1'b0;
      out_sig_25_sv2v_reg <= 1'b0;
      out_sig_24_sv2v_reg <= 1'b0;
      out_sig_23_sv2v_reg <= 1'b0;
      out_sig_22_sv2v_reg <= 1'b0;
      out_sig_21_sv2v_reg <= 1'b0;
      out_sig_20_sv2v_reg <= 1'b0;
      out_sig_19_sv2v_reg <= 1'b0;
      out_sig_18_sv2v_reg <= 1'b0;
      out_sig_17_sv2v_reg <= 1'b0;
      out_sig_16_sv2v_reg <= 1'b0;
      out_sig_15_sv2v_reg <= 1'b0;
      out_sig_14_sv2v_reg <= 1'b0;
      out_sig_13_sv2v_reg <= 1'b0;
      out_sig_12_sv2v_reg <= 1'b0;
      out_sig_11_sv2v_reg <= 1'b0;
      out_sig_10_sv2v_reg <= 1'b0;
      out_sig_9_sv2v_reg <= 1'b0;
      out_sig_8_sv2v_reg <= 1'b0;
      out_sig_7_sv2v_reg <= 1'b0;
      out_sig_6_sv2v_reg <= 1'b0;
      out_sig_5_sv2v_reg <= 1'b0;
      out_sig_4_sv2v_reg <= 1'b0;
      out_sig_3_sv2v_reg <= 1'b0;
      out_sig_2_sv2v_reg <= 1'b0;
      out_sig_1_sv2v_reg <= 1'b0;
    end else if(N297) begin
      out_sig_0_sv2v_reg <= N298;
      out_sig_26_sv2v_reg <= N357;
      out_sig_25_sv2v_reg <= N358;
      out_sig_24_sv2v_reg <= N359;
      out_sig_23_sv2v_reg <= N353;
      out_sig_22_sv2v_reg <= N352;
      out_sig_21_sv2v_reg <= N351;
      out_sig_20_sv2v_reg <= N350;
      out_sig_19_sv2v_reg <= N349;
      out_sig_18_sv2v_reg <= N348;
      out_sig_17_sv2v_reg <= N347;
      out_sig_16_sv2v_reg <= N346;
      out_sig_15_sv2v_reg <= N345;
      out_sig_14_sv2v_reg <= N344;
      out_sig_13_sv2v_reg <= N343;
      out_sig_12_sv2v_reg <= N342;
      out_sig_11_sv2v_reg <= N341;
      out_sig_10_sv2v_reg <= N340;
      out_sig_9_sv2v_reg <= N339;
      out_sig_8_sv2v_reg <= N338;
      out_sig_7_sv2v_reg <= N337;
      out_sig_6_sv2v_reg <= N336;
      out_sig_5_sv2v_reg <= N335;
      out_sig_4_sv2v_reg <= N334;
      out_sig_3_sv2v_reg <= N333;
      out_sig_2_sv2v_reg <= N332;
      out_sig_1_sv2v_reg <= N331;
    end 
    if(N59) begin
      rem_Z_25_sv2v_reg <= 1'b0;
      rem_Z_24_sv2v_reg <= 1'b0;
      rem_Z_23_sv2v_reg <= 1'b0;
      rem_Z_22_sv2v_reg <= 1'b0;
      rem_Z_21_sv2v_reg <= 1'b0;
      rem_Z_20_sv2v_reg <= 1'b0;
      rem_Z_19_sv2v_reg <= 1'b0;
      rem_Z_18_sv2v_reg <= 1'b0;
      rem_Z_17_sv2v_reg <= 1'b0;
      rem_Z_16_sv2v_reg <= 1'b0;
      rem_Z_15_sv2v_reg <= 1'b0;
      rem_Z_14_sv2v_reg <= 1'b0;
      rem_Z_13_sv2v_reg <= 1'b0;
      rem_Z_12_sv2v_reg <= 1'b0;
      rem_Z_11_sv2v_reg <= 1'b0;
      rem_Z_10_sv2v_reg <= 1'b0;
      rem_Z_9_sv2v_reg <= 1'b0;
      rem_Z_8_sv2v_reg <= 1'b0;
      rem_Z_7_sv2v_reg <= 1'b0;
      rem_Z_6_sv2v_reg <= 1'b0;
      rem_Z_5_sv2v_reg <= 1'b0;
      rem_Z_4_sv2v_reg <= 1'b0;
      rem_Z_3_sv2v_reg <= 1'b0;
      rem_Z_2_sv2v_reg <= 1'b0;
      rem_Z_1_sv2v_reg <= 1'b0;
      rem_Z_0_sv2v_reg <= 1'b0;
    end else if(N269) begin
      rem_Z_25_sv2v_reg <= N296;
      rem_Z_24_sv2v_reg <= N295;
      rem_Z_23_sv2v_reg <= N294;
      rem_Z_22_sv2v_reg <= N293;
      rem_Z_21_sv2v_reg <= N292;
      rem_Z_20_sv2v_reg <= N291;
      rem_Z_19_sv2v_reg <= N290;
      rem_Z_18_sv2v_reg <= N289;
      rem_Z_17_sv2v_reg <= N288;
      rem_Z_16_sv2v_reg <= N287;
      rem_Z_15_sv2v_reg <= N286;
      rem_Z_14_sv2v_reg <= N285;
      rem_Z_13_sv2v_reg <= N284;
      rem_Z_12_sv2v_reg <= N283;
      rem_Z_11_sv2v_reg <= N282;
      rem_Z_10_sv2v_reg <= N281;
      rem_Z_9_sv2v_reg <= N280;
      rem_Z_8_sv2v_reg <= N279;
      rem_Z_7_sv2v_reg <= N278;
      rem_Z_6_sv2v_reg <= N277;
      rem_Z_5_sv2v_reg <= N276;
      rem_Z_4_sv2v_reg <= N275;
      rem_Z_3_sv2v_reg <= N274;
      rem_Z_2_sv2v_reg <= N273;
      rem_Z_1_sv2v_reg <= N272;
      rem_Z_0_sv2v_reg <= N271;
    end 
  end


endmodule



module roundRawFNToRecFN_expWidth8_sigWidth24_options0
(
  control,
  invalidExc,
  infiniteExc,
  in_isNaN,
  in_isInf,
  in_isZero,
  in_sign,
  in_sExp,
  in_sig,
  roundingMode,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [9:0] in_sExp;
  input [26:0] in_sig;
  input [2:0] roundingMode;
  output [32:0] out;
  output [4:0] exceptionFlags;
  input invalidExc;
  input infiniteExc;
  input in_isNaN;
  input in_isInf;
  input in_isZero;
  input in_sign;
  wire [32:0] out;
  wire [4:0] exceptionFlags;

  roundAnyRawFNToRecFN_inExpWidth8_inSigWidth26_outExpWidth8_outSigWidth24_options0
  roundAnyRawFNToRecFN
  (
    .control(control[0]),
    .invalidExc(invalidExc),
    .infiniteExc(infiniteExc),
    .in_isNaN(in_isNaN),
    .in_isInf(in_isInf),
    .in_isZero(in_isZero),
    .in_sign(in_sign),
    .in_sExp(in_sExp),
    .in_sig(in_sig),
    .roundingMode(roundingMode),
    .out(out),
    .exceptionFlags(exceptionFlags)
  );


endmodule



module divSqrtRecFN_small_expWidth8_sigWidth24
(
  nReset,
  clock,
  control,
  inReady,
  inValid,
  sqrtOp,
  a,
  b,
  roundingMode,
  outValid,
  sqrtOpOut,
  out,
  exceptionFlags
);

  input [0:0] control;
  input [32:0] a;
  input [32:0] b;
  input [2:0] roundingMode;
  output [32:0] out;
  output [4:0] exceptionFlags;
  input nReset;
  input clock;
  input inValid;
  input sqrtOp;
  output inReady;
  output outValid;
  output sqrtOpOut;
  wire [32:0] out;
  wire [4:0] exceptionFlags;
  wire inReady,outValid,sqrtOpOut,invalidExc,infiniteExc,out_isNaN,out_isInf,
  out_isZero,out_sign;
  wire [2:0] roundingModeOut;
  wire [9:0] out_sExp;
  wire [26:0] out_sig;

  divSqrtRecFNToRaw_small_expWidth8_sigWidth24_options0
  divSqrtRecFNToRaw
  (
    .nReset(nReset),
    .clock(clock),
    .control(control[0]),
    .inReady(inReady),
    .inValid(inValid),
    .sqrtOp(sqrtOp),
    .a(a),
    .b(b),
    .roundingMode(roundingMode),
    .outValid(outValid),
    .sqrtOpOut(sqrtOpOut),
    .roundingModeOut(roundingModeOut),
    .invalidExc(invalidExc),
    .infiniteExc(infiniteExc),
    .out_isNaN(out_isNaN),
    .out_isInf(out_isInf),
    .out_isZero(out_isZero),
    .out_sign(out_sign),
    .out_sExp(out_sExp),
    .out_sig(out_sig)
  );


  roundRawFNToRecFN_expWidth8_sigWidth24_options0
  roundRawOut
  (
    .control(control[0]),
    .invalidExc(invalidExc),
    .infiniteExc(infiniteExc),
    .in_isNaN(out_isNaN),
    .in_isInf(out_isInf),
    .in_isZero(out_isZero),
    .in_sign(out_sign),
    .in_sExp(out_sExp),
    .in_sig(out_sig),
    .roundingMode(roundingModeOut),
    .out(out),
    .exceptionFlags(exceptionFlags)
  );


endmodule



module fpu_fdiv_fsqrt
(
  clk_i,
  reset_i,
  v_i,
  rd_i,
  rm_i,
  fp_rs1_i,
  fp_rs2_i,
  fsqrt_i,
  ready_o,
  v_o,
  result_o,
  rd_o,
  yumi_i,
  fflags_o_invalid_,
  fflags_o_div_zero_,
  fflags_o_overflow_,
  fflags_o_underflow_,
  fflags_o_inexact_
);

  input [4:0] rd_i;
  input [2:0] rm_i;
  input [32:0] fp_rs1_i;
  input [32:0] fp_rs2_i;
  output [32:0] result_o;
  output [4:0] rd_o;
  input clk_i;
  input reset_i;
  input v_i;
  input fsqrt_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output fflags_o_invalid_;
  output fflags_o_div_zero_;
  output fflags_o_overflow_;
  output fflags_o_underflow_;
  output fflags_o_inexact_;
  wire [32:0] result_o;
  wire [4:0] rd_o;
  wire ready_o,v_o,fflags_o_invalid_,fflags_o_div_zero_,fflags_o_overflow_,
  fflags_o_underflow_,fflags_o_inexact_,N0,N1,N2,N3,N4,N5,N6,_0_net_,ready_lo,v_li,v_lo,N7,N8,
  N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,
  N29;
  wire [1:0] ds_state_n,ds_state_r;
  reg rd_o_4_sv2v_reg,rd_o_3_sv2v_reg,rd_o_2_sv2v_reg,rd_o_1_sv2v_reg,rd_o_0_sv2v_reg,
  ds_state_r_1_sv2v_reg,ds_state_r_0_sv2v_reg;
  assign rd_o[4] = rd_o_4_sv2v_reg;
  assign rd_o[3] = rd_o_3_sv2v_reg;
  assign rd_o[2] = rd_o_2_sv2v_reg;
  assign rd_o[1] = rd_o_1_sv2v_reg;
  assign rd_o[0] = rd_o_0_sv2v_reg;
  assign ds_state_r[1] = ds_state_r_1_sv2v_reg;
  assign ds_state_r[0] = ds_state_r_0_sv2v_reg;

  divSqrtRecFN_small_expWidth8_sigWidth24
  ds0
  (
    .nReset(_0_net_),
    .clock(clk_i),
    .control(1'b1),
    .inReady(ready_lo),
    .inValid(v_li),
    .sqrtOp(fsqrt_i),
    .a(fp_rs1_i),
    .b(fp_rs2_i),
    .roundingMode(rm_i),
    .outValid(v_lo),
    .out(result_o),
    .exceptionFlags({ fflags_o_invalid_, fflags_o_div_zero_, fflags_o_overflow_, fflags_o_underflow_, fflags_o_inexact_ })
  );

  assign N9 = N7 & N8;
  assign N10 = ds_state_r[1] | N8;
  assign N12 = N7 | ds_state_r[0];
  assign N14 = ds_state_r[1] & ds_state_r[0];
  assign { N21, N20, N19, N18, N17 } = (N0)? rd_i : 
                                       (N16)? rd_o : 1'b0;
  assign N0 = N15;
  assign { N25, N24 } = (N1)? { N26, 1'b0 } : 
                        (N2)? ds_state_r : 1'b0;
  assign N1 = v_lo;
  assign N2 = N23;
  assign ready_o = (N3)? ready_lo : 
                   (N4)? 1'b0 : 
                   (N5)? 1'b0 : 
                   (N6)? 1'b0 : 1'b0;
  assign N3 = N9;
  assign N4 = N11;
  assign N5 = N13;
  assign N6 = N14;
  assign v_li = (N3)? v_i : 
                (N4)? 1'b0 : 
                (N5)? 1'b0 : 
                (N6)? 1'b0 : 1'b0;
  assign ds_state_n = (N3)? { 1'b0, N22 } : 
                      (N4)? { N25, N24 } : 
                      (N5)? { N26, 1'b0 } : 
                      (N6)? { 1'b0, 1'b0 } : 1'b0;
  assign v_o = (N3)? 1'b0 : 
               (N4)? v_lo : 
               (N5)? 1'b1 : 
               (N6)? 1'b0 : 1'b0;
  assign _0_net_ = ~reset_i;
  assign N7 = ~ds_state_r[1];
  assign N8 = ~ds_state_r[0];
  assign N11 = ~N10;
  assign N13 = ~N12;
  assign N15 = ready_lo & v_i;
  assign N16 = ~N15;
  assign N22 = ready_lo & v_i;
  assign N23 = ~v_lo;
  assign N26 = ~yumi_i;
  assign N27 = N11 | N13;
  assign N28 = N27 | N14;
  assign N29 = ~N28;

  always @(posedge clk_i) begin
    if(reset_i) begin
      rd_o_4_sv2v_reg <= 1'b0;
      rd_o_3_sv2v_reg <= 1'b0;
      rd_o_2_sv2v_reg <= 1'b0;
      rd_o_1_sv2v_reg <= 1'b0;
      rd_o_0_sv2v_reg <= 1'b0;
    end else if(N29) begin
      rd_o_4_sv2v_reg <= N21;
      rd_o_3_sv2v_reg <= N20;
      rd_o_2_sv2v_reg <= N19;
      rd_o_1_sv2v_reg <= N18;
      rd_o_0_sv2v_reg <= N17;
    end 
    if(reset_i) begin
      ds_state_r_1_sv2v_reg <= 1'b0;
      ds_state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      ds_state_r_1_sv2v_reg <= ds_state_n[1];
      ds_state_r_0_sv2v_reg <= ds_state_n[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p44
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [43:0] data_i;
  output [43:0] data_o;
  input clk_i;
  input reset_i;
  wire [43:0] data_o;
  reg data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,
  data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,
  data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_43_sv2v_reg <= 1'b0;
      data_o_42_sv2v_reg <= 1'b0;
      data_o_41_sv2v_reg <= 1'b0;
      data_o_40_sv2v_reg <= 1'b0;
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_width_p32
(
  clk_i,
  data_i,
  data_o
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  wire [31:0] data_o;
  reg data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p1024_data_width_p32_latch_last_read_p1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [9:0] addr_i;
  input [31:0] data_i;
  input [3:0] write_mask_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [31:0] data_o;

//  fakeram130_1024x32 fakeram1
//(
//   data_o,
//   addr_i,
//   w_i,
//   data_i,
//   write_mask_i,
//   clk_i,
//   vi_i);

  hard_mem_1rw_byte_mask_d1024_w32_wrapper
  \macro.mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_reset_width_p1
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p32_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input en_i;
  wire [31:0] data_o;
  reg data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,
  data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,
  data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p32
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input en_i;
  wire [31:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p32_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_dff_reset_width_p40
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [39:0] data_i;
  output [39:0] data_o;
  input clk_i;
  input reset_i;
  wire [39:0] data_o;
  reg data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_39_sv2v_reg <= 1'b0;
      data_o_38_sv2v_reg <= 1'b0;
      data_o_37_sv2v_reg <= 1'b0;
      data_o_36_sv2v_reg <= 1'b0;
      data_o_35_sv2v_reg <= 1'b0;
      data_o_34_sv2v_reg <= 1'b0;
      data_o_33_sv2v_reg <= 1'b0;
      data_o_32_sv2v_reg <= 1'b0;
      data_o_31_sv2v_reg <= 1'b0;
      data_o_30_sv2v_reg <= 1'b0;
      data_o_29_sv2v_reg <= 1'b0;
      data_o_28_sv2v_reg <= 1'b0;
      data_o_27_sv2v_reg <= 1'b0;
      data_o_26_sv2v_reg <= 1'b0;
      data_o_25_sv2v_reg <= 1'b0;
      data_o_24_sv2v_reg <= 1'b0;
      data_o_23_sv2v_reg <= 1'b0;
      data_o_22_sv2v_reg <= 1'b0;
      data_o_21_sv2v_reg <= 1'b0;
      data_o_20_sv2v_reg <= 1'b0;
      data_o_19_sv2v_reg <= 1'b0;
      data_o_18_sv2v_reg <= 1'b0;
      data_o_17_sv2v_reg <= 1'b0;
      data_o_16_sv2v_reg <= 1'b0;
      data_o_15_sv2v_reg <= 1'b0;
      data_o_14_sv2v_reg <= 1'b0;
      data_o_13_sv2v_reg <= 1'b0;
      data_o_12_sv2v_reg <= 1'b0;
      data_o_11_sv2v_reg <= 1'b0;
      data_o_10_sv2v_reg <= 1'b0;
      data_o_9_sv2v_reg <= 1'b0;
      data_o_8_sv2v_reg <= 1'b0;
      data_o_7_sv2v_reg <= 1'b0;
      data_o_6_sv2v_reg <= 1'b0;
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_reset_width_p6
(
  clk_i,
  reset_i,
  data_i,
  data_o
);

  input [5:0] data_i;
  output [5:0] data_o;
  input clk_i;
  input reset_i;
  wire [5:0] data_o;
  reg data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_o_5_sv2v_reg <= 1'b0;
      data_o_4_sv2v_reg <= 1'b0;
      data_o_3_sv2v_reg <= 1'b0;
      data_o_2_sv2v_reg <= 1'b0;
      data_o_1_sv2v_reg <= 1'b0;
      data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_mux_width_p32_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[63] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[62] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[61] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[60] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[59] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[58] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[57] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[56] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[55] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[54] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[53] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[52] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[51] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[50] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[49] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[48] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[47] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[46] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[45] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[44] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[43] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[42] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[41] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[40] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[39] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[38] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[37] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[36] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[35] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[34] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[33] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[32] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_scan_width_p3_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [2:0] i;
  output [2:0] o;
  wire [2:0] o;
  wire t_1__2_,t_1__1_,t_1__0_;
  assign t_1__2_ = i[0] | 1'b0;
  assign t_1__1_ = i[1] | i[0];
  assign t_1__0_ = i[2] | i[1];
  assign o[0] = t_1__2_ | 1'b0;
  assign o[1] = t_1__1_ | 1'b0;
  assign o[2] = t_1__0_ | t_1__2_;

endmodule



module bsg_priority_encode_one_hot_out_width_p3_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [2:0] i;
  output [2:0] o;
  output v_o;
  wire [2:0] o;
  wire v_o,N0,N1;
  wire [1:1] scan_lo;

  bsg_scan_width_p3_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo[1:1], o[0:0] })
  );

  assign o[2] = v_o & N0;
  assign N0 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N1;
  assign N1 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p3_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [2:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o;
  wire v_o,v_1__0_;
  assign v_1__0_ = i[1] | i[0];
  assign addr_o[1] = 1'b0 | i[2];
  assign v_o = addr_o[1] | v_1__0_;
  assign addr_o[0] = i[1] | 1'b0;

endmodule



module bsg_priority_encode_width_p3_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [2:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o;
  wire v_o;
  wire [2:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p3_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p3_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module vanilla_core_data_width_p32_dmem_size_p1024_icache_entries_p1024_icache_tag_width_p12_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_credit_counter_width_p6_fwd_fifo_els_p3
(
  clk_i,
  reset_i,
  pc_init_val_i,
  remote_req_o,
  remote_req_v_o,
  remote_req_credit_i,
  icache_v_i,
  icache_pc_i,
  icache_instr_i,
  icache_yumi_o,
  ifetch_v_i,
  ifetch_instr_i,
  remote_dmem_v_i,
  remote_dmem_w_i,
  remote_dmem_addr_i,
  remote_dmem_mask_i,
  remote_dmem_data_i,
  remote_dmem_data_o,
  remote_dmem_yumi_o,
  float_remote_load_resp_rd_i,
  float_remote_load_resp_data_i,
  float_remote_load_resp_v_i,
  float_remote_load_resp_force_i,
  float_remote_load_resp_yumi_o,
  int_remote_load_resp_rd_i,
  int_remote_load_resp_data_i,
  int_remote_load_resp_v_i,
  int_remote_load_resp_force_i,
  int_remote_load_resp_yumi_o,
  invalid_eva_access_i,
  remote_interrupt_set_i,
  remote_interrupt_clear_i,
  remote_interrupt_pending_bit_o,
  out_credits_used_i,
  cfg_pod_x_o,
  cfg_pod_y_o,
  global_x_i,
  global_y_i
);

  input [21:0] pc_init_val_i;
  output [83:0] remote_req_o;
  input [21:0] icache_pc_i;
  input [31:0] icache_instr_i;
  input [31:0] ifetch_instr_i;
  input [9:0] remote_dmem_addr_i;
  input [3:0] remote_dmem_mask_i;
  input [31:0] remote_dmem_data_i;
  output [31:0] remote_dmem_data_o;
  input [4:0] float_remote_load_resp_rd_i;
  input [31:0] float_remote_load_resp_data_i;
  input [4:0] int_remote_load_resp_rd_i;
  input [31:0] int_remote_load_resp_data_i;
  input [5:0] out_credits_used_i;
  output [2:0] cfg_pod_x_o;
  output [3:0] cfg_pod_y_o;
  input [6:0] global_x_i;
  input [6:0] global_y_i;
  input clk_i;
  input reset_i;
  input remote_req_credit_i;
  input icache_v_i;
  input ifetch_v_i;
  input remote_dmem_v_i;
  input remote_dmem_w_i;
  input float_remote_load_resp_v_i;
  input float_remote_load_resp_force_i;
  input int_remote_load_resp_v_i;
  input int_remote_load_resp_force_i;
  input invalid_eva_access_i;
  input remote_interrupt_set_i;
  input remote_interrupt_clear_i;
  output remote_req_v_o;
  output icache_yumi_o;
  output remote_dmem_yumi_o;
  output float_remote_load_resp_yumi_o;
  output int_remote_load_resp_yumi_o;
  output remote_interrupt_pending_bit_o;
  wire [83:0] remote_req_o;
  wire [31:0] remote_dmem_data_o,icache_winstr,instruction,mcsr_data_lo,mem_addr_op2,fsw_data,
  rs1_forward_val,wb_data_r,mem_result,exe_result,rs2_forward_val,rs1_val_to_exe,
  rs2_val_to_exe,alu_result,alu_or_csr_result,idiv_result_lo,lsu_dmem_data_lo,
  lsu_mem_addr_sent_lo,imul_result_lo,fpu_int_result_lo,mem_data_n,mem_data_r,
  dmem_data_li,local_load_data_r,local_load_packed_data,wb_data_n,flw_wb_data_n,
  flw_wb_data_r,flw_data;
  wire [2:0] cfg_pod_x_o,float_rf_read,frm_r,has_forward_data_rs1,has_forward_data_rs2,
  fpu_rm;
  wire [3:0] cfg_pod_y_o,lsu_dmem_mask_lo,dmem_mask_li;
  wire remote_req_v_o,icache_yumi_o,remote_dmem_yumi_o,float_remote_load_resp_yumi_o,
  int_remote_load_resp_yumi_o,remote_interrupt_pending_bit_o,N0,N1,N2,N3,N4,N5,N6,
  N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,icache_v_li,icache_w_li,
  icache_flush,icache_miss,icache_flush_r_lo,int_sb_score,int_sb_clear,int_dependency,
  float_rf_wen,float_sb_score,float_sb_clear,float_dependency,fcsr_v_li,fcsr_data_v_lo,
  fcsr_fflags_li_1__invalid_,fcsr_fflags_li_1__div_zero_,
  fcsr_fflags_li_1__overflow_,fcsr_fflags_li_1__underflow_,fcsr_fflags_li_1__inexact_,mcsr_we_li,
  mcsr_instr_executed_li,mcsr_interrupt_entered_li,mcsr_mret_called_li,mstatus_r_mpie_,
  mstatus_r_mie_,mip_r_trace_,mie_r_trace_,mie_r_remote_,remote_interrupt_ready,
  trace_interrupt_ready,interrupt_ready,is_amo_or_lr_op,N40,N41,N42,N43,aq_r,aq_set,
  aq_clear,N44,N45,N46,N47,N48,N49,frs1_forward_v,frs2_forward_v,frs3_forward_v,
  rs1_forward_v,N50,rs2_forward_v,N51,N52,N53,N54,N55,alu_jump_now,
  jalr_prediction_write_en,N56,N57,idiv_v_li,idiv_ready_lo,idiv_v_lo,idiv_yumi_li,lsu_remote_req_v_lo,
  lsu_dmem_v_lo,lsu_dmem_w_lo,lsu_reserve_lo,npc_write_en,branch_under_predict,
  branch_over_predict,branch_mispredict,N58,jalr_mispredict,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,stall_fpu2_li,imul_v_lo,fpu_float_v_lo,
  fpu_float_fflags_lo_invalid_,fpu_float_fflags_lo_div_zero_,fpu_float_fflags_lo_overflow_,
  fpu_float_fflags_lo_underflow_,fpu_float_fflags_lo_inexact_,fpu1_v_r,
  fpu_int_fflags_lo_invalid_,fpu_int_fflags_lo_div_zero_,fpu_int_fflags_lo_overflow_,
  fpu_int_fflags_lo_underflow_,fpu_int_fflags_lo_inexact_,fdiv_fsqrt_v_li,fdiv_fsqrt_ready_lo,
  fdiv_fsqrt_v_lo,fdiv_fsqrt_fflags_lo_invalid_,fdiv_fsqrt_fflags_lo_div_zero_,
  fdiv_fsqrt_fflags_lo_overflow_,fdiv_fsqrt_fflags_lo_underflow_,fdiv_fsqrt_fflags_lo_inexact_,
  fdiv_fsqrt_yumi_li,dmem_v_li,dmem_w_li,local_load_en,local_load_en_r,reserved_r,
  make_reserve,break_reserve,N70,N71,N72,N73,N74,N75,select_remote_flw,
  stall_depend_long_op,stall_depend_local_load,stall_depend_imul,stall_bypass,stall_lr_aq,
  stall_fence,stall_amo_aq,stall_amo_rl,stall_remote_req,stall_remote_credit,
  stall_fdiv_busy,stall_idiv_busy,stall_fcsr,stall_id,stall_icache_store,
  stall_remote_ld_wb,stall_ifetch_wait,stall_remote_flw_wb,stall_all,flush,icache_miss_in_pipe,
  reset_r,reset_down,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,read_icache,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,rf_read_en,
  local_load_in_exe,int_remote_load_in_exe,float_remote_load_in_exe,fdiv_fsqrt_in_fp_exe,
  id_rs1_equal_exe_rd,id_rs2_equal_exe_rd,id_rs3_equal_exe_rd,
  id_rs1_equal_fp_exe_rd,id_rs2_equal_fp_exe_rd,id_rs3_equal_fp_exe_rd,id_rs1_equal_mem_rd,
  id_rs2_equal_mem_rd,id_rs3_equal_mem_rd,id_rs1_equal_wb_rd,id_rs2_equal_wb_rd,N152,
  rs1_sb_clear_now,N153,frs2_sb_clear_now,N154,N155,N156,N157,N158,stall_bypass_fp_frs,
  N159,stall_bypass_fp_rs1,N160,N161,N162,stall_bypass_int_frs2,N163,
  local_mem_op_restore,id_remote_req_op,memory_op_issued,N164,N165,N166,N167,N168,N169,N170,N171,
  N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,
  N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,
  N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,
  N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,
  N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,
  N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,
  N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,
  N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,
  N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,
  N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,
  N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,
  N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,
  N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,
  N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,
  N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,
  N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,
  N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,
  N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,
  N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,
  N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,
  N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,
  N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,mem_result_valid,N519,
  N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,
  N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,
  N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,
  N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
  N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,
  N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,
  N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,
  N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,
  N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,
  N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,
  N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,
  N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,
  N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,
  N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
  N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,
  N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,
  N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,
  N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,
  N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,
  N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,
  N840,N841,N842,N843,N844,N845,N846;
  wire [21:0] icache_w_pc,pc_n,jalr_prediction,pred_or_jump_addr,pc_r,pc_plus4,mepc_r,
  alu_jalr_addr,npc_n,npc_r;
  wire [30:0] decode;
  wire [10:0] fp_decode;
  wire [139:0] id_n,id_r;
  wire [1:0] int_rf_read,fcsr_fflags_v_li,rs1_forward_sel,rs2_forward_sel,
  remote_req_counter_r,remote_req_available;
  wire [63:0] int_rf_rdata;
  wire [4:0] float_rf_waddr,float_sb_score_id,float_sb_clear_id,aq_rd_r,idiv_rd_lo,
  imul_rd_lo,fpu_float_rd_lo,fpu1_rd_r,fdiv_fsqrt_rd_lo;
  wire [32:0] float_rf_wdata,frs1_select_val,frs1_to_fp_exe,frs2_to_fp_exe,frs3_to_fp_exe,
  fpu_float_result_lo,fdiv_fsqrt_result_lo,flw_recoded_data;
  wire [98:0] float_rf_rdata,fp_exe_data_n,fp_exe_data_r;
  wire [7:0] fcsr_data_lo;
  wire [5:0] credit_limit_r,flw_wb_ctrl_n,flw_wb_ctrl_r;
  wire [224:0] exe_r,exe_n;
  wire [43:0] mem_ctrl_r,mem_ctrl_n;
  wire [39:0] wb_ctrl_r,wb_ctrl_n;
  wire [9:0] lsu_dmem_addr_lo,dmem_addr_li,reserved_addr_r;
  wire [18:0] fp_exe_ctrl_n,fp_exe_ctrl_r;
  reg aq_rd_r_4_sv2v_reg,aq_rd_r_3_sv2v_reg,aq_rd_r_2_sv2v_reg,aq_rd_r_1_sv2v_reg,
  aq_rd_r_0_sv2v_reg,aq_r_sv2v_reg,reserved_addr_r_9_sv2v_reg,
  reserved_addr_r_8_sv2v_reg,reserved_addr_r_7_sv2v_reg,reserved_addr_r_6_sv2v_reg,
  reserved_addr_r_5_sv2v_reg,reserved_addr_r_4_sv2v_reg,reserved_addr_r_3_sv2v_reg,
  reserved_addr_r_2_sv2v_reg,reserved_addr_r_1_sv2v_reg,reserved_addr_r_0_sv2v_reg,reserved_r_sv2v_reg,
  remote_req_counter_r_1_sv2v_reg,remote_req_counter_r_0_sv2v_reg;
  assign aq_rd_r[4] = aq_rd_r_4_sv2v_reg;
  assign aq_rd_r[3] = aq_rd_r_3_sv2v_reg;
  assign aq_rd_r[2] = aq_rd_r_2_sv2v_reg;
  assign aq_rd_r[1] = aq_rd_r_1_sv2v_reg;
  assign aq_rd_r[0] = aq_rd_r_0_sv2v_reg;
  assign aq_r = aq_r_sv2v_reg;
  assign reserved_addr_r[9] = reserved_addr_r_9_sv2v_reg;
  assign reserved_addr_r[8] = reserved_addr_r_8_sv2v_reg;
  assign reserved_addr_r[7] = reserved_addr_r_7_sv2v_reg;
  assign reserved_addr_r[6] = reserved_addr_r_6_sv2v_reg;
  assign reserved_addr_r[5] = reserved_addr_r_5_sv2v_reg;
  assign reserved_addr_r[4] = reserved_addr_r_4_sv2v_reg;
  assign reserved_addr_r[3] = reserved_addr_r_3_sv2v_reg;
  assign reserved_addr_r[2] = reserved_addr_r_2_sv2v_reg;
  assign reserved_addr_r[1] = reserved_addr_r_1_sv2v_reg;
  assign reserved_addr_r[0] = reserved_addr_r_0_sv2v_reg;
  assign reserved_r = reserved_r_sv2v_reg;
  assign remote_req_counter_r[1] = remote_req_counter_r_1_sv2v_reg;
  assign remote_req_counter_r[0] = remote_req_counter_r_0_sv2v_reg;

  icache_icache_tag_width_p12_icache_entries_p1024
  icache0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(icache_v_li),
    .w_i(icache_w_li),
    .flush_i(icache_flush),
    .w_pc_i(icache_w_pc),
    .w_instr_i(icache_winstr),
    .pc_i(pc_n),
    .jalr_prediction_i(jalr_prediction),
    .instr_o(instruction),
    .pred_or_jump_addr_o(pred_or_jump_addr),
    .pc_r_o(pc_r),
    .icache_miss_o(icache_miss),
    .icache_flush_r_o(icache_flush_r_lo)
  );


  cl_decode
  decode0
  (
    .instruction_i(instruction),
    .decode_o(decode),
    .fp_decode_o(fp_decode)
  );


  bsg_dff_reset_width_p140
  id_pipeline
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(id_n),
    .data_o(id_r)
  );


  regfile_width_p32_els_p32_num_rs_p2_x0_tied_to_zero_p1
  int_rf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(wb_ctrl_r[39]),
    .w_addr_i(wb_ctrl_r[38:34]),
    .w_data_i(wb_data_r),
    .r_v_i(int_rf_read),
    .r_addr_i(instruction[24:15]),
    .r_data_o(int_rf_rdata)
  );


  scoreboard_els_p32_num_src_port_p2_num_clear_port_p1_x0_tied_to_zero_p1
  int_sb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .src_id_i(id_r[68:59]),
    .dest_id_i(id_r[55:51]),
    .op_reads_rf_i({ id_r[42:42], id_r[43:43] }),
    .op_writes_rf_i(id_r[41]),
    .score_i(int_sb_score),
    .score_id_i(exe_r[140:136]),
    .clear_i(int_sb_clear),
    .clear_id_i(wb_ctrl_r[38:34]),
    .dependency_o(int_dependency)
  );


  regfile_width_p33_els_p32_num_rs_p3_x0_tied_to_zero_p0
  float_rf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(float_rf_wen),
    .w_addr_i(float_rf_waddr),
    .w_data_i(float_rf_wdata),
    .r_v_i(float_rf_read),
    .r_addr_i({ instruction[31:27], instruction[24:15] }),
    .r_data_o(float_rf_rdata)
  );


  scoreboard_els_p32_num_src_port_p3_num_clear_port_p1_x0_tied_to_zero_p0
  float_sb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .src_id_i({ id_r[75:71], id_r[68:59] }),
    .dest_id_i(id_r[55:51]),
    .op_reads_rf_i({ id_r[17:17], id_r[18:18], id_r[19:19] }),
    .op_writes_rf_i(id_r[16]),
    .score_i(float_sb_score),
    .score_id_i(float_sb_score_id),
    .clear_i(float_sb_clear),
    .clear_id_i(float_sb_clear_id),
    .dependency_o(float_dependency)
  );


  fcsr
  fcsr0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(fcsr_v_li),
    .funct3_i(id_r[58:56]),
    .rs1_i(id_r[63:59]),
    .data_i(rs1_val_to_exe[7:0]),
    .addr_i(id_r[75:64]),
    .data_o(fcsr_data_lo),
    .data_v_o(fcsr_data_v_lo),
    .fflags_v_i(fcsr_fflags_v_li),
    .fflags_i({ fcsr_fflags_li_1__invalid_, fcsr_fflags_li_1__div_zero_, fcsr_fflags_li_1__overflow_, fcsr_fflags_li_1__underflow_, fcsr_fflags_li_1__inexact_, fpu_int_fflags_lo_invalid_, fpu_int_fflags_lo_div_zero_, fpu_int_fflags_lo_overflow_, fpu_int_fflags_lo_underflow_, fpu_int_fflags_lo_inexact_ }),
    .frm_o(frm_r)
  );


  mcsr_pc_width_p22_credit_counter_width_p6_cfg_pod_width_p7
  mcsr0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .remote_interrupt_set_i(remote_interrupt_set_i),
    .remote_interrupt_clear_i(remote_interrupt_clear_i),
    .we_i(mcsr_we_li),
    .addr_i(id_r[75:64]),
    .funct3_i(id_r[58:56]),
    .data_i(rs1_val_to_exe),
    .rs1_i(id_r[63:59]),
    .data_o(mcsr_data_lo),
    .cfg_pod_reset_val_i({ global_y_i[6:3], global_x_i[6:4] }),
    .cfg_pod_r_o({ cfg_pod_y_o, cfg_pod_x_o }),
    .instr_executed_i(mcsr_instr_executed_li),
    .interrupt_entered_i(mcsr_interrupt_entered_li),
    .mret_called_i(mcsr_mret_called_li),
    .npc_r_i(npc_r),
    .mepc_r_o(mepc_r),
    .credit_limit_o(credit_limit_r),
    .mstatus_r_o_mpie_(mstatus_r_mpie_),
    .mstatus_r_o_mie_(mstatus_r_mie_),
    .mip_r_o_trace_(mip_r_trace_),
    .mip_r_o_remote_(remote_interrupt_pending_bit_o),
    .mie_r_o_trace_(mie_r_trace_),
    .mie_r_o_remote_(mie_r_remote_)
  );


  bsg_mux_width_p33_els_p2
  frs1_select_mux
  (
    .data_i({ 1'b0, int_rf_rdata[31:0], float_rf_rdata[32:0] }),
    .sel_i(id_r[43]),
    .data_o(frs1_select_val)
  );


  bsg_mux_width_p33_els_p2
  frs1_fwd_mux
  (
    .data_i({ float_rf_wdata, frs1_select_val }),
    .sel_i(frs1_forward_v),
    .data_o(frs1_to_fp_exe)
  );


  bsg_mux_width_p33_els_p2
  frs2_fwd_mux
  (
    .data_i({ float_rf_wdata, float_rf_rdata[65:33] }),
    .sel_i(frs2_forward_v),
    .data_o(frs2_to_fp_exe)
  );


  bsg_mux_width_p33_els_p2
  frs3_fwd_mux
  (
    .data_i({ float_rf_wdata, float_rf_rdata[98:66] }),
    .sel_i(frs3_forward_v),
    .data_o(frs3_to_fp_exe)
  );


  recFNToFN_expWidth8_sigWidth24
  frs2_to_fn
  (
    .in(float_rf_rdata[65:33]),
    .out(fsw_data)
  );


  bsg_mux_width_p32_els_p3
  exe_rs1_fwd_mux
  (
    .data_i({ wb_data_r, mem_result, exe_result }),
    .sel_i(rs1_forward_sel),
    .data_o(rs1_forward_val)
  );


  bsg_mux_width_p32_els_p3
  exe_rs2_fwd_mux
  (
    .data_i({ wb_data_r, mem_result, exe_result }),
    .sel_i(rs2_forward_sel),
    .data_o(rs2_forward_val)
  );


  bsg_dff_reset_width_p225
  exe_pipeline
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(exe_n),
    .data_o(exe_r)
  );


  alu_pc_width_p22
  alu0
  (
    .rs1_i(exe_r[97:66]),
    .rs2_i(exe_r[65:34]),
    .pc_plus4_i(exe_r[224:193]),
    .op_i(exe_r[160:129]),
    .result_o(alu_result),
    .jalr_addr_o(alu_jalr_addr),
    .jump_now_o(alu_jump_now)
  );


  bsg_dff_reset_en_bypass_width_p22
  jalr_pred_dff
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(jalr_prediction_write_en),
    .data_i(exe_r[216:195]),
    .data_o(jalr_prediction)
  );


  idiv
  idiv0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(idiv_v_li),
    .rs1_i(exe_r[97:66]),
    .rs2_i(exe_r[65:34]),
    .rd_i(exe_r[140:136]),
    .op_i(exe_r[115:114]),
    .ready_o(idiv_ready_lo),
    .v_o(idiv_v_lo),
    .rd_o(idiv_rd_lo),
    .result_o(idiv_result_lo),
    .yumi_i(idiv_yumi_li)
  );


  lsu_data_width_p32_pc_width_p22_dmem_size_p1024
  lsu0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .exe_decode_i(exe_r[128:98]),
    .exe_rs1_i(exe_r[97:66]),
    .exe_rs2_i(exe_r[65:34]),
    .exe_rd_i(exe_r[140:136]),
    .mem_offset_i(exe_r[33:2]),
    .pc_plus4_i(exe_r[224:193]),
    .icache_miss_i(exe_r[1]),
    .remote_req_o(remote_req_o),
    .remote_req_v_o(lsu_remote_req_v_lo),
    .dmem_v_o(lsu_dmem_v_lo),
    .dmem_w_o(lsu_dmem_w_lo),
    .dmem_addr_o(lsu_dmem_addr_lo),
    .dmem_data_o(lsu_dmem_data_lo),
    .dmem_mask_o(lsu_dmem_mask_lo),
    .reserve_o(lsu_reserve_lo),
    .mem_addr_sent_o(lsu_mem_addr_sent_lo)
  );


  bsg_dff_en_bypass_width_p22
  npc_dff
  (
    .clk_i(clk_i),
    .en_i(npc_write_en),
    .data_i(npc_n),
    .data_o(npc_r)
  );

  assign N58 = alu_jalr_addr != exe_r[184:163];

  bsg_dff_reset_width_p19
  fp_exe_ctrl_pipeline
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(fp_exe_ctrl_n),
    .data_o(fp_exe_ctrl_r)
  );


  bsg_dff_width_p99
  fp_exe_data_pipeline
  (
    .clk_i(clk_i),
    .data_i(fp_exe_data_n),
    .data_o(fp_exe_data_r)
  );


  fpu_float
  fpu_float0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .stall_fpu1_i(stall_all),
    .stall_fpu2_i(stall_fpu2_li),
    .imul_v_i(exe_r[117]),
    .imul_rs1_i(exe_r[97:66]),
    .imul_rs2_i(exe_r[65:34]),
    .imul_rd_i(exe_r[140:136]),
    .fp_v_i(fp_exe_ctrl_r[13]),
    .fpu_float_op_i(fp_exe_ctrl_r[9:6]),
    .fp_rs1_i(fp_exe_data_r[98:66]),
    .fp_rs2_i(fp_exe_data_r[65:33]),
    .fp_rs3_i(fp_exe_data_r[32:0]),
    .fp_rd_i(fp_exe_ctrl_r[18:14]),
    .fp_rm_i(fp_exe_ctrl_r[2:0]),
    .imul_v_o(imul_v_lo),
    .imul_result_o(imul_result_lo),
    .imul_rd_o(imul_rd_lo),
    .fp_v_o(fpu_float_v_lo),
    .fp_result_o(fpu_float_result_lo),
    .fp_rd_o(fpu_float_rd_lo),
    .fpu1_v_r_o(fpu1_v_r),
    .fpu1_rd_o(fpu1_rd_r),
    .fp_fflags_o_invalid_(fpu_float_fflags_lo_invalid_),
    .fp_fflags_o_div_zero_(fpu_float_fflags_lo_div_zero_),
    .fp_fflags_o_overflow_(fpu_float_fflags_lo_overflow_),
    .fp_fflags_o_underflow_(fpu_float_fflags_lo_underflow_),
    .fp_fflags_o_inexact_(fpu_float_fflags_lo_inexact_)
  );


  fpu_int
  fpu_int0
  (
    .fp_rs1_i(fp_exe_data_r[98:66]),
    .fp_rs2_i(fp_exe_data_r[65:33]),
    .fpu_int_op_i(fp_exe_ctrl_r[5:3]),
    .fp_rm_i(fp_exe_ctrl_r[2:0]),
    .result_o(fpu_int_result_lo),
    .fflags_o_invalid_(fpu_int_fflags_lo_invalid_),
    .fflags_o_div_zero_(fpu_int_fflags_lo_div_zero_),
    .fflags_o_overflow_(fpu_int_fflags_lo_overflow_),
    .fflags_o_underflow_(fpu_int_fflags_lo_underflow_),
    .fflags_o_inexact_(fpu_int_fflags_lo_inexact_)
  );


  fpu_fdiv_fsqrt
  fpu_fdiv_fsqrt0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(fdiv_fsqrt_v_li),
    .rd_i(fp_exe_ctrl_r[18:14]),
    .rm_i(fp_exe_ctrl_r[2:0]),
    .fp_rs1_i(fp_exe_data_r[98:66]),
    .fp_rs2_i(fp_exe_data_r[65:33]),
    .fsqrt_i(fp_exe_ctrl_r[10]),
    .ready_o(fdiv_fsqrt_ready_lo),
    .v_o(fdiv_fsqrt_v_lo),
    .result_o(fdiv_fsqrt_result_lo),
    .rd_o(fdiv_fsqrt_rd_lo),
    .yumi_i(fdiv_fsqrt_yumi_li),
    .fflags_o_invalid_(fdiv_fsqrt_fflags_lo_invalid_),
    .fflags_o_div_zero_(fdiv_fsqrt_fflags_lo_div_zero_),
    .fflags_o_overflow_(fdiv_fsqrt_fflags_lo_overflow_),
    .fflags_o_underflow_(fdiv_fsqrt_fflags_lo_underflow_),
    .fflags_o_inexact_(fdiv_fsqrt_fflags_lo_inexact_)
  );


  bsg_dff_reset_width_p44
  mem_ctrl_pipeline
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(mem_ctrl_n),
    .data_o(mem_ctrl_r)
  );


  bsg_dff_width_p32
  mem_data_pipeline
  (
    .clk_i(clk_i),
    .data_i(mem_data_n),
    .data_o(mem_data_r)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p1024_data_width_p32_latch_last_read_p1
  dmem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(dmem_v_li),
    .w_i(dmem_w_li),
    .addr_i(dmem_addr_li),
    .data_i(dmem_data_li),
    .write_mask_i(dmem_mask_li),
    .data_o(remote_dmem_data_o)
  );


  bsg_dff_reset_width_p1
  local_load_en_dff
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(local_load_en),
    .data_o(local_load_en_r)
  );


  bsg_dff_en_bypass_width_p32
  local_load_buffer
  (
    .clk_i(clk_i),
    .en_i(local_load_en_r),
    .data_i(remote_dmem_data_o),
    .data_o(local_load_data_r)
  );


  load_packer
  local_lp
  (
    .mem_data_i(local_load_data_r),
    .unsigned_load_i(mem_ctrl_r[34]),
    .byte_load_i(mem_ctrl_r[36]),
    .hex_load_i(mem_ctrl_r[35]),
    .part_sel_i(mem_ctrl_r[2:1]),
    .load_data_o(local_load_packed_data)
  );


  bsg_dff_reset_width_p40
  wb_ctrl_pipeline
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(wb_ctrl_n),
    .data_o(wb_ctrl_r)
  );


  bsg_dff_width_p32
  wb_data_pipeline
  (
    .clk_i(clk_i),
    .data_i(wb_data_n),
    .data_o(wb_data_r)
  );


  bsg_dff_reset_width_p6
  flw_wb_ctrl_pipeline
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(flw_wb_ctrl_n),
    .data_o(flw_wb_ctrl_r)
  );


  bsg_dff_width_p32
  flw_wb_data_pipeline
  (
    .clk_i(clk_i),
    .data_i(flw_wb_data_n),
    .data_o(flw_wb_data_r)
  );


  bsg_mux_width_p32_els_p2
  flw_recFN_mux
  (
    .data_i({ float_remote_load_resp_data_i, flw_wb_data_r }),
    .sel_i(select_remote_flw),
    .data_o(flw_data)
  );


  fNToRecFN_expWidth8_sigWidth24
  flw_to_RecFN
  (
    .in(flw_data),
    .out(flw_recoded_data)
  );


  bsg_dff_width_p1
  reset_dff
  (
    .clk_i(clk_i),
    .data_i(reset_i),
    .data_o(reset_r)
  );

  assign id_rs1_equal_exe_rd = id_r[63:59] == exe_r[140:136];
  assign id_rs2_equal_exe_rd = id_r[68:64] == exe_r[140:136];
  assign id_rs3_equal_exe_rd = id_r[75:71] == exe_r[140:136];
  assign id_rs1_equal_fp_exe_rd = id_r[63:59] == fp_exe_ctrl_r[18:14];
  assign id_rs2_equal_fp_exe_rd = id_r[68:64] == fp_exe_ctrl_r[18:14];
  assign id_rs3_equal_fp_exe_rd = id_r[75:71] == fp_exe_ctrl_r[18:14];
  assign id_rs1_equal_mem_rd = id_r[63:59] == mem_ctrl_r[43:39];
  assign id_rs2_equal_mem_rd = id_r[68:64] == mem_ctrl_r[43:39];
  assign id_rs3_equal_mem_rd = id_r[75:71] == mem_ctrl_r[43:39];
  assign id_rs1_equal_wb_rd = id_r[63:59] == wb_ctrl_r[38:34];
  assign id_rs2_equal_wb_rd = id_r[68:64] == wb_ctrl_r[38:34];
  assign N152 = id_r[63:59] == wb_ctrl_r[38:34];
  assign N153 = id_r[68:64] == float_sb_clear_id;
  assign N156 = id_r[63:59] == fpu1_rd_r;
  assign N157 = id_r[68:64] == fpu1_rd_r;
  assign N158 = id_r[75:71] == fpu1_rd_r;
  assign N159 = id_r[63:59] == imul_rd_lo;
  assign N160 = id_r[68:64] == fpu1_rd_r;
  assign N161 = id_r[68:64] == fpu_float_rd_lo;
  assign N162 = id_r[68:64] == flw_wb_ctrl_r[4:0];
  assign N171 = remote_req_available == 1'b0;
  assign N178 = { N177, N176, N175, N174, N173, N172 } >= credit_limit_r;
  assign N184 = id_r[63:59] == float_rf_waddr;
  assign N185 = id_r[68:64] == float_rf_waddr;
  assign N186 = id_r[75:71] == float_rf_waddr;
  assign N187 = imul_rd_lo == id_r[63:59];

  bsg_priority_encode_width_p3_lo_to_hi_p1
  rs1_forward_pe0
  (
    .i(has_forward_data_rs1),
    .addr_o(rs1_forward_sel),
    .v_o(rs1_forward_v)
  );

  assign N188 = imul_rd_lo == id_r[68:64];

  bsg_priority_encode_width_p3_lo_to_hi_p1
  rs2_forward_pe0
  (
    .i(has_forward_data_rs2),
    .addr_o(rs2_forward_sel),
    .v_o(rs2_forward_v)
  );

  assign N189 = wb_ctrl_r[38:34] == aq_rd_r;
  assign N514 = reserved_addr_r == dmem_addr_li;
  assign N597 = ~exe_r[136];
  assign N598 = exe_r[139] | exe_r[140];
  assign N599 = exe_r[138] | N598;
  assign N600 = exe_r[137] | N599;
  assign N601 = N597 | N600;
  assign N602 = ~N601;
  assign N603 = ~exe_r[138];
  assign N604 = ~exe_r[136];
  assign N605 = exe_r[139] | exe_r[140];
  assign N606 = N603 | N605;
  assign N607 = exe_r[137] | N606;
  assign N608 = N604 | N607;
  assign N609 = ~N608;
  assign N610 = id_r[57] & id_r[58];
  assign N611 = id_r[56] & N610;
  assign N612 = id_r[67] | id_r[68];
  assign N613 = id_r[66] | N612;
  assign N614 = id_r[65] | N613;
  assign N615 = id_r[64] | N614;
  assign N616 = out_credits_used_i[4] | out_credits_used_i[5];
  assign N617 = out_credits_used_i[3] | N616;
  assign N618 = out_credits_used_i[2] | N617;
  assign N619 = out_credits_used_i[1] | N618;
  assign N620 = out_credits_used_i[0] | N619;
  assign N621 = ~id_r[64];
  assign N622 = id_r[74] | id_r[75];
  assign N623 = id_r[73] | N622;
  assign N624 = id_r[72] | N623;
  assign N625 = id_r[71] | N624;
  assign N626 = id_r[70] | N625;
  assign N627 = id_r[69] | N626;
  assign N628 = id_r[68] | N627;
  assign N629 = id_r[67] | N628;
  assign N630 = id_r[66] | N629;
  assign N631 = id_r[65] | N630;
  assign N632 = N621 | N631;
  assign N633 = ~N632;
  assign N634 = ~id_r[65];
  assign N635 = ~id_r[64];
  assign N636 = id_r[74] | id_r[75];
  assign N637 = id_r[73] | N636;
  assign N638 = id_r[72] | N637;
  assign N639 = id_r[71] | N638;
  assign N640 = id_r[70] | N639;
  assign N641 = id_r[69] | N640;
  assign N642 = id_r[68] | N641;
  assign N643 = id_r[67] | N642;
  assign N644 = id_r[66] | N643;
  assign N645 = N634 | N644;
  assign N646 = N635 | N645;
  assign N647 = ~N646;
  assign N648 = id_r[62] | id_r[63];
  assign N649 = id_r[61] | N648;
  assign N650 = id_r[60] | N649;
  assign N651 = id_r[59] | N650;
  assign { N177, N176, N175, N174, N173, N172 } = out_credits_used_i + lsu_remote_req_v_lo;
  assign { N165, N164 } = remote_req_counter_r + remote_req_credit_i;
  assign pc_plus4 = pc_r + 1'b1;
  assign { N167, N166 } = { N165, N164 } + local_mem_op_restore;
  assign remote_req_available = { N167, N166 } + invalid_eva_access_i;
  assign { N170, N169 } = remote_req_available - memory_op_issued;
  assign mem_addr_op2 = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                        (N43)? { id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:69], id_r[55:51] } : 
                        (N41)? { id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:75], id_r[75:64] } : 1'b0;
  assign N0 = is_amo_or_lr_op;
  assign N46 = (N1)? 1'b1 : 
               (N49)? 1'b1 : 
               (N45)? 1'b0 : 1'b0;
  assign N1 = aq_set;
  assign N47 = (N1)? 1'b1 : 
               (N49)? 1'b0 : 
               (N45)? 1'b0 : 1'b0;
  assign rs1_val_to_exe = (N2)? rs1_forward_val : 
                          (N3)? int_rf_rdata[31:0] : 1'b0;
  assign N2 = rs1_forward_v;
  assign N3 = N50;
  assign rs2_val_to_exe = (N4)? fsw_data : 
                          (N55)? rs2_forward_val : 
                          (N53)? int_rf_rdata[63:32] : 1'b0;
  assign N4 = N51;
  assign alu_or_csr_result = (N5)? exe_r[65:34] : 
                             (N57)? alu_result : 1'b0;
  assign N5 = N56;
  assign npc_n = (N6)? alu_jalr_addr : 
                 (N66)? mepc_r : 
                 (N69)? exe_r[184:163] : 
                 (N64)? exe_r[216:195] : 1'b0;
  assign N6 = N60;
  assign N72 = (N7)? 1'b1 : 
               (N75)? 1'b1 : 
               (N71)? 1'b0 : 1'b0;
  assign N7 = make_reserve;
  assign N73 = (N7)? 1'b1 : 
               (N75)? 1'b0 : 
               (N71)? 1'b0 : 1'b0;
  assign { N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88 } = (N8)? exe_r[184:163] : 
                                                                                                                                      (N9)? exe_r[216:195] : 1'b0;
  assign N8 = alu_jump_now;
  assign N9 = N661;
  assign pc_n = (N10)? pc_init_val_i : 
                (N111)? wb_ctrl_r[24:3] : 
                (N114)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N87 } : 
                (N117)? mepc_r : 
                (N120)? { N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88 } : 
                (N123)? alu_jalr_addr : 
                (N126)? pred_or_jump_addr : 
                (N129)? pred_or_jump_addr : 
                (N86)? pc_plus4 : 1'b0;
  assign N10 = reset_down;
  assign read_icache = (N11)? wb_ctrl_r[33] : 
                       (N131)? 1'b1 : 1'b0;
  assign N11 = N130;
  assign icache_w_pc = (N12)? mem_ctrl_r[24:3] : 
                       (N13)? icache_pc_i : 1'b0;
  assign N12 = ifetch_v_i;
  assign N13 = N132;
  assign icache_winstr = (N12)? ifetch_instr_i : 
                         (N13)? icache_instr_i : 1'b0;
  assign id_n = (N14)? id_r : 
                (N142)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N145)? id_r : 
                (N148)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N151)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, pc_plus4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N140)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, pc_plus4, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, pred_or_jump_addr, 1'b0, 1'b0, instruction, decode, fp_decode, 1'b0, 1'b1 } : 1'b0;
  assign N14 = N135;
  assign N155 = (N15)? rs1_sb_clear_now : 
                (N154)? frs2_sb_clear_now : 1'b0;
  assign N15 = id_r[20];
  assign stall_bypass = (N15)? N163 : 
                        (N154)? stall_bypass_int_frs2 : 1'b0;
  assign N181 = (N16)? N180 : 
                (N17)? 1'b1 : 1'b0;
  assign N16 = fdiv_fsqrt_ready_lo;
  assign N17 = N179;
  assign N183 = (N18)? exe_r[116] : 
                (N19)? 1'b1 : 1'b0;
  assign N18 = idiv_ready_lo;
  assign N19 = N182;
  assign { N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198 } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fcsr_data_lo } : 
                                                                                                                                                                                                              (N21)? mcsr_data_lo : 1'b0;
  assign N20 = fcsr_data_v_lo;
  assign N21 = N197;
  assign { N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230 } = (N22)? { N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198 } : 
                                                                                                                                                                                                              (N196)? rs2_val_to_exe : 1'b0;
  assign N22 = id_r[15];
  assign { N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262 } = (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N488)? { id_r[139:108], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, id_r[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N195)? { id_r[139:13], rs1_val_to_exe, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, mem_addr_op2, id_r[1:0] } : 1'b0;
  assign N23 = N193;
  assign exe_n = (N24)? exe_r : 
                 (N25)? { N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262 } : 1'b0;
  assign N24 = N191;
  assign N25 = N190;
  assign npc_write_en = (N24)? 1'b0 : 
                        (N25)? N192 : 1'b0;
  assign exe_result = (N26)? fpu_int_result_lo : 
                      (N489)? alu_or_csr_result : 1'b0;
  assign N26 = fp_exe_ctrl_r[12];
  assign fpu_rm = (N27)? frm_r : 
                  (N490)? id_r[58:56] : 1'b0;
  assign N27 = N611;
  assign { fp_exe_ctrl_n[18:14], fp_exe_ctrl_n[9:0] } = (N494)? { id_r[55:51], id_r[8:2], fpu_rm } : 
                                                        (N495)? { fp_exe_ctrl_r[18:14], fp_exe_ctrl_r[9:0] } : 1'b0;
  assign fp_exe_ctrl_n[13:10] = (N28)? fp_exe_ctrl_r[13:10] : 
                                (N497)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N494)? id_r[12:9] : 1'b0;
  assign N28 = N492;
  assign fp_exe_data_n = (N28)? fp_exe_data_r : 
                         (N497)? fp_exe_data_r : 
                         (N494)? { frs1_to_fp_exe, frs2_to_fp_exe, frs3_to_fp_exe } : 1'b0;
  assign float_sb_score_id = (N29)? fp_exe_ctrl_r[18:14] : 
                             (N30)? exe_r[140:136] : 1'b0;
  assign N29 = fdiv_fsqrt_in_fp_exe;
  assign N30 = N498;
  assign mem_ctrl_n = (N31)? mem_ctrl_r : 
                      (N505)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N508)? { fp_exe_ctrl_r[18:14], 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N503)? { exe_r[140:136], exe_r[126:126], exe_r[101:101], exe_r[123:121], local_load_in_exe, lsu_mem_addr_sent_lo, exe_r[1:1] } : 1'b0;
  assign N31 = N500;
  assign mem_data_n = (N31)? mem_data_r : 
                      (N505)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N508)? fpu_int_result_lo : 
                      (N503)? alu_or_csr_result : 1'b0;
  assign fcsr_fflags_v_li[0] = (N31)? 1'b0 : 
                               (N505)? 1'b0 : 
                               (N508)? 1'b1 : 
                               (N503)? 1'b0 : 1'b0;
  assign dmem_v_li = (N32)? remote_dmem_v_i : 
                     (N513)? 1'b1 : 
                     (N511)? remote_dmem_v_i : 1'b0;
  assign N32 = N509;
  assign dmem_w_li = (N32)? remote_dmem_w_i : 
                     (N513)? lsu_dmem_w_lo : 
                     (N511)? remote_dmem_w_i : 1'b0;
  assign dmem_addr_li = (N32)? remote_dmem_addr_i : 
                        (N513)? lsu_dmem_addr_lo : 
                        (N511)? remote_dmem_addr_i : 1'b0;
  assign dmem_data_li = (N32)? remote_dmem_data_i : 
                        (N513)? lsu_dmem_data_lo : 
                        (N511)? remote_dmem_data_i : 1'b0;
  assign dmem_mask_li = (N32)? remote_dmem_mask_i : 
                        (N513)? lsu_dmem_mask_lo : 
                        (N511)? remote_dmem_mask_i : 1'b0;
  assign remote_dmem_yumi_o = (N32)? remote_dmem_v_i : 
                              (N513)? 1'b0 : 
                              (N511)? remote_dmem_v_i : 1'b0;
  assign local_load_en = (N32)? 1'b0 : 
                         (N513)? N692 : 
                         (N511)? 1'b0 : 1'b0;
  assign mem_result = (N33)? imul_result_lo : 
                      (N518)? local_load_packed_data : 
                      (N516)? mem_data_r : 1'b0;
  assign N33 = imul_v_lo;
  assign { N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528 } = (N34)? local_load_packed_data : 
                                                                                                                                                                                                              (N527)? mem_data_r : 1'b0;
  assign N34 = mem_ctrl_r[33];
  assign { wb_ctrl_n[39:34], wb_ctrl_n[0:0] } = (N35)? { 1'b1, int_remote_load_resp_rd_i, 1'b1 } : 
                                                (wb_ctrl_n[33])? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N566)? { 1'b1, imul_rd_lo, 1'b0 } : 
                                                (N568)? { 1'b1, mem_ctrl_r[43:39], 1'b0 } : 
                                                (N571)? { 1'b1, int_remote_load_resp_rd_i, 1'b1 } : 
                                                (N574)? { 1'b1, idiv_rd_lo, 1'b1 } : 
                                                (N525)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N35 = int_remote_load_resp_force_i;
  assign wb_ctrl_n[32:1] = (wb_ctrl_n[33])? mem_ctrl_r[32:1] : 
                           (N561)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign wb_data_n = (N35)? int_remote_load_resp_data_i : 
                     (wb_ctrl_n[33])? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N566)? imul_result_lo : 
                     (N568)? { N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528 } : 
                     (N571)? int_remote_load_resp_data_i : 
                     (N574)? idiv_result_lo : 
                     (N525)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stall_remote_ld_wb = (N35)? N526 : 
                              (N562)? 1'b0 : 
                              (N36)? 1'b0 : 
                              (N36)? 1'b0 : 
                              (N36)? 1'b0 : 
                              (N36)? 1'b0 : 
                              (N36)? 1'b0 : 1'b0;
  assign N36 = 1'b0;
  assign int_remote_load_resp_yumi_o = (N35)? 1'b1 : 
                                       (wb_ctrl_n[33])? 1'b0 : 
                                       (N566)? 1'b0 : 
                                       (N568)? 1'b0 : 
                                       (N571)? 1'b1 : 
                                       (N563)? 1'b0 : 
                                       (N36)? 1'b0 : 1'b0;
  assign idiv_yumi_li = (N35)? 1'b0 : 
                        (wb_ctrl_n[33])? 1'b0 : 
                        (N566)? 1'b0 : 
                        (N568)? 1'b0 : 
                        (N571)? 1'b0 : 
                        (N574)? 1'b1 : 
                        (N525)? 1'b0 : 1'b0;
  assign flw_wb_ctrl_n = (N37)? flw_wb_ctrl_r : 
                         (N38)? { mem_ctrl_r[37:37], mem_ctrl_r[43:39] } : 1'b0;
  assign N37 = N576;
  assign N38 = N575;
  assign flw_wb_data_n = (N37)? flw_wb_data_r : 
                         (N38)? local_load_data_r : 1'b0;
  assign select_remote_flw = (N39)? 1'b1 : 
                             (N587)? 1'b0 : 
                             (N590)? 1'b0 : 
                             (N593)? 1'b0 : 
                             (N596)? 1'b1 : 
                             (N581)? 1'b0 : 1'b0;
  assign N39 = float_remote_load_resp_force_i;
  assign float_rf_wen = (N39)? 1'b1 : 
                        (N587)? 1'b1 : 
                        (N590)? 1'b1 : 
                        (N593)? 1'b1 : 
                        (N596)? 1'b1 : 
                        (N581)? 1'b0 : 1'b0;
  assign float_rf_waddr = (N39)? float_remote_load_resp_rd_i : 
                          (N587)? flw_wb_ctrl_r[4:0] : 
                          (N590)? fpu_float_rd_lo : 
                          (N593)? fdiv_fsqrt_rd_lo : 
                          (N596)? float_remote_load_resp_rd_i : 
                          (N581)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign float_rf_wdata = (N39)? flw_recoded_data : 
                          (N587)? flw_recoded_data : 
                          (N590)? fpu_float_result_lo : 
                          (N593)? fdiv_fsqrt_result_lo : 
                          (N596)? flw_recoded_data : 
                          (N581)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign float_remote_load_resp_yumi_o = (N39)? 1'b1 : 
                                         (N587)? 1'b0 : 
                                         (N590)? 1'b0 : 
                                         (N593)? 1'b0 : 
                                         (N596)? 1'b1 : 
                                         (N581)? 1'b0 : 1'b0;
  assign stall_remote_flw_wb = (N39)? N582 : 
                               (N583)? 1'b0 : 
                               (N36)? 1'b0 : 
                               (N36)? 1'b0 : 
                               (N36)? 1'b0 : 
                               (N36)? 1'b0 : 1'b0;
  assign float_sb_clear = (N39)? 1'b1 : 
                          (N587)? 1'b0 : 
                          (N590)? 1'b0 : 
                          (N593)? 1'b1 : 
                          (N596)? 1'b1 : 
                          (N581)? 1'b0 : 1'b0;
  assign float_sb_clear_id = (N593)? fdiv_fsqrt_rd_lo : 
                             (N585)? float_remote_load_resp_rd_i : 1'b0;
  assign fcsr_fflags_v_li[1] = (N39)? 1'b0 : 
                               (N587)? 1'b0 : 
                               (N590)? 1'b1 : 
                               (N593)? 1'b1 : 
                               (N586)? 1'b0 : 
                               (N36)? 1'b0 : 1'b0;
  assign { fcsr_fflags_li_1__invalid_, fcsr_fflags_li_1__div_zero_, fcsr_fflags_li_1__overflow_, fcsr_fflags_li_1__underflow_, fcsr_fflags_li_1__inexact_ } = (N39)? { fpu_float_fflags_lo_invalid_, fpu_float_fflags_lo_div_zero_, fpu_float_fflags_lo_overflow_, fpu_float_fflags_lo_underflow_, fpu_float_fflags_lo_inexact_ } : 
                                                                                                                                                              (N587)? { fpu_float_fflags_lo_invalid_, fpu_float_fflags_lo_div_zero_, fpu_float_fflags_lo_overflow_, fpu_float_fflags_lo_underflow_, fpu_float_fflags_lo_inexact_ } : 
                                                                                                                                                              (N590)? { fpu_float_fflags_lo_invalid_, fpu_float_fflags_lo_div_zero_, fpu_float_fflags_lo_overflow_, fpu_float_fflags_lo_underflow_, fpu_float_fflags_lo_inexact_ } : 
                                                                                                                                                              (N593)? { fdiv_fsqrt_fflags_lo_invalid_, fdiv_fsqrt_fflags_lo_div_zero_, fdiv_fsqrt_fflags_lo_overflow_, fdiv_fsqrt_fflags_lo_underflow_, fdiv_fsqrt_fflags_lo_inexact_ } : 
                                                                                                                                                              (N586)? { fpu_float_fflags_lo_invalid_, fpu_float_fflags_lo_div_zero_, fpu_float_fflags_lo_overflow_, fpu_float_fflags_lo_underflow_, fpu_float_fflags_lo_inexact_ } : 
                                                                                                                                                              (N36)? { fpu_float_fflags_lo_invalid_, fpu_float_fflags_lo_div_zero_, fpu_float_fflags_lo_overflow_, fpu_float_fflags_lo_underflow_, fpu_float_fflags_lo_inexact_ } : 1'b0;
  assign fdiv_fsqrt_yumi_li = (N39)? 1'b0 : 
                              (N587)? 1'b0 : 
                              (N590)? 1'b0 : 
                              (N593)? 1'b1 : 
                              (N586)? 1'b0 : 
                              (N36)? 1'b0 : 1'b0;
  assign remote_interrupt_ready = remote_interrupt_pending_bit_o & mie_r_remote_;
  assign trace_interrupt_ready = mip_r_trace_ & mie_r_trace_;
  assign interrupt_ready = N653 & N656;
  assign N653 = mstatus_r_mie_ & N652;
  assign N652 = remote_interrupt_ready | trace_interrupt_ready;
  assign N656 = ~N655;
  assign N655 = N654 | wb_ctrl_r[33];
  assign N654 = exe_r[1] | mem_ctrl_r[0];
  assign is_amo_or_lr_op = N657 | id_r[25];
  assign N657 = id_r[26] | id_r[27];
  assign N40 = id_r[39] | is_amo_or_lr_op;
  assign N41 = ~N40;
  assign N42 = ~is_amo_or_lr_op;
  assign N43 = id_r[39] & N42;
  assign N44 = aq_clear | aq_set;
  assign N45 = ~N44;
  assign N48 = ~aq_set;
  assign N49 = aq_clear & N48;
  assign N50 = ~rs1_forward_v;
  assign N51 = id_r[18];
  assign N52 = rs2_forward_v | N51;
  assign N53 = ~N52;
  assign N54 = ~N51;
  assign N55 = rs2_forward_v & N54;
  assign jalr_prediction_write_en = N658 & N659;
  assign N658 = exe_r[119] | exe_r[118];
  assign N659 = N602 | N609;
  assign N56 = exe_r[100];
  assign N57 = ~N56;
  assign branch_under_predict = alu_jump_now & N660;
  assign N660 = ~exe_r[129];
  assign branch_over_predict = N661 & exe_r[129];
  assign N661 = ~alu_jump_now;
  assign branch_mispredict = N662 & exe_r[120];
  assign N662 = branch_under_predict | branch_over_predict;
  assign jalr_mispredict = exe_r[118] & N58;
  assign N59 = exe_r[119] | N663;
  assign N663 = exe_r[120] & alu_jump_now;
  assign N60 = exe_r[118];
  assign N61 = exe_r[99];
  assign N62 = N61 | N60;
  assign N63 = N59 | N62;
  assign N64 = ~N63;
  assign N65 = ~N60;
  assign N66 = N61 & N65;
  assign N67 = ~N61;
  assign N68 = N65 & N67;
  assign N69 = N59 & N68;
  assign N70 = break_reserve | make_reserve;
  assign N71 = ~N70;
  assign N74 = ~make_reserve;
  assign N75 = break_reserve & N74;
  assign stall_id = N674 | stall_fcsr;
  assign N674 = N673 | stall_idiv_busy;
  assign N673 = N672 | stall_fdiv_busy;
  assign N672 = N671 | stall_remote_credit;
  assign N671 = N670 | stall_remote_req;
  assign N670 = N669 | stall_amo_rl;
  assign N669 = N668 | stall_amo_aq;
  assign N668 = N667 | stall_fence;
  assign N667 = N666 | stall_lr_aq;
  assign N666 = N665 | stall_bypass;
  assign N665 = N664 | stall_depend_imul;
  assign N664 = stall_depend_long_op | stall_depend_local_load;
  assign stall_all = N678 | stall_remote_flw_wb;
  assign N678 = N677 | 1'b0;
  assign N677 = N676 | stall_ifetch_wait;
  assign N676 = N675 | stall_remote_ld_wb;
  assign N675 = stall_icache_store | 1'b0;
  assign flush = N680 | interrupt_ready;
  assign N680 = N679 | exe_r[99];
  assign N679 = branch_mispredict | jalr_mispredict;
  assign icache_miss_in_pipe = N682 | wb_ctrl_r[33];
  assign N682 = N681 | mem_ctrl_r[0];
  assign N681 = id_r[1] | exe_r[1];
  assign reset_down = reset_r & N683;
  assign N683 = ~reset_i;
  assign N76 = decode[22] & instruction[0];
  assign N77 = decode[21] | decode[20];
  assign N78 = exe_r[99];
  assign N79 = wb_ctrl_r[33] | reset_down;
  assign N80 = interrupt_ready | N79;
  assign N81 = N78 | N80;
  assign N82 = branch_mispredict | N81;
  assign N83 = jalr_mispredict | N82;
  assign N84 = N76 | N83;
  assign N85 = N77 | N84;
  assign N86 = ~N85;
  assign N87 = ~remote_interrupt_ready;
  assign N110 = ~reset_down;
  assign N111 = wb_ctrl_r[33] & N110;
  assign N112 = ~wb_ctrl_r[33];
  assign N113 = N110 & N112;
  assign N114 = interrupt_ready & N113;
  assign N115 = ~interrupt_ready;
  assign N116 = N113 & N115;
  assign N117 = N78 & N116;
  assign N118 = ~N78;
  assign N119 = N116 & N118;
  assign N120 = branch_mispredict & N119;
  assign N121 = ~branch_mispredict;
  assign N122 = N119 & N121;
  assign N123 = jalr_mispredict & N122;
  assign N124 = ~jalr_mispredict;
  assign N125 = N122 & N124;
  assign N126 = N76 & N125;
  assign N127 = ~N76;
  assign N128 = N125 & N127;
  assign N129 = N77 & N128;
  assign N130 = icache_miss_in_pipe & N684;
  assign N684 = ~flush;
  assign N131 = ~N130;
  assign icache_v_li = N685 | N690;
  assign N685 = icache_v_i | ifetch_v_i;
  assign N690 = N687 & N689;
  assign N687 = read_icache & N686;
  assign N686 = ~stall_all;
  assign N689 = ~N688;
  assign N688 = stall_id & N684;
  assign icache_w_li = icache_v_i | ifetch_v_i;
  assign N132 = ~ifetch_v_i;
  assign icache_yumi_o = icache_v_i & N132;
  assign icache_flush = flush | icache_miss_in_pipe;
  assign stall_icache_store = icache_v_i & icache_yumi_o;
  assign N133 = reset_down | flush;
  assign N134 = icache_miss_in_pipe | icache_flush_r_lo;
  assign N135 = stall_all;
  assign N136 = N133 | N135;
  assign N137 = stall_id | N136;
  assign N138 = N134 | N137;
  assign N139 = icache_miss | N138;
  assign N140 = ~N139;
  assign N141 = ~N135;
  assign N142 = N133 & N141;
  assign N143 = ~N133;
  assign N144 = N141 & N143;
  assign N145 = stall_id & N144;
  assign N146 = ~stall_id;
  assign N147 = N144 & N146;
  assign N148 = N134 & N147;
  assign N149 = ~N134;
  assign N150 = N147 & N149;
  assign N151 = icache_miss & N150;
  assign rf_read_en = ~N691;
  assign N691 = stall_id | stall_all;
  assign int_rf_read[0] = id_n[43] & rf_read_en;
  assign int_rf_read[1] = id_n[42] & rf_read_en;
  assign float_rf_read[0] = id_n[19] & rf_read_en;
  assign float_rf_read[1] = id_n[18] & rf_read_en;
  assign float_rf_read[2] = id_n[17] & rf_read_en;
  assign local_load_in_exe = lsu_dmem_v_lo & N692;
  assign N692 = ~lsu_dmem_w_lo;
  assign int_remote_load_in_exe = N693 & exe_r[126];
  assign N693 = lsu_remote_req_v_lo & exe_r[125];
  assign float_remote_load_in_exe = N694 & exe_r[101];
  assign N694 = lsu_remote_req_v_lo & exe_r[125];
  assign fdiv_fsqrt_in_fp_exe = fp_exe_ctrl_r[11] | fp_exe_ctrl_r[10];
  assign rs1_sb_clear_now = N696 & N651;
  assign N696 = N695 & int_sb_clear;
  assign N695 = id_r[43] & N152;
  assign frs2_sb_clear_now = N697 & float_sb_clear;
  assign N697 = id_r[18] & N153;
  assign N154 = ~id_r[20];
  assign stall_depend_long_op = N698 | N155;
  assign N698 = int_dependency | float_dependency;
  assign stall_depend_local_load = local_load_in_exe & N714;
  assign N714 = N711 | N713;
  assign N711 = N708 | N710;
  assign N708 = N705 | N707;
  assign N705 = N701 | N704;
  assign N701 = N700 & N651;
  assign N700 = N699 & exe_r[126];
  assign N699 = id_r[43] & id_rs1_equal_exe_rd;
  assign N704 = N703 & N615;
  assign N703 = N702 & exe_r[126];
  assign N702 = id_r[42] & id_rs2_equal_exe_rd;
  assign N707 = N706 & exe_r[101];
  assign N706 = id_r[19] & id_rs1_equal_exe_rd;
  assign N710 = N709 & exe_r[101];
  assign N709 = id_r[18] & id_rs2_equal_exe_rd;
  assign N713 = N712 & exe_r[101];
  assign N712 = id_r[17] & id_rs3_equal_exe_rd;
  assign stall_depend_imul = exe_r[117] & N719;
  assign N719 = N716 | N718;
  assign N716 = N715 & N651;
  assign N715 = id_r[43] & id_rs1_equal_exe_rd;
  assign N718 = N717 & N615;
  assign N717 = id_r[42] & id_rs2_equal_exe_rd;
  assign stall_bypass_fp_frs = N742 | N744;
  assign N742 = N739 | N741;
  assign N739 = N736 | N738;
  assign N736 = N733 | N735;
  assign N733 = N730 | N732;
  assign N730 = N727 | N729;
  assign N727 = N724 | N726;
  assign N724 = N721 | N723;
  assign N721 = N720 & fp_exe_ctrl_r[13];
  assign N720 = id_r[19] & id_rs1_equal_fp_exe_rd;
  assign N723 = N722 & fp_exe_ctrl_r[13];
  assign N722 = id_r[18] & id_rs2_equal_fp_exe_rd;
  assign N726 = N725 & fp_exe_ctrl_r[13];
  assign N725 = id_r[17] & id_rs3_equal_fp_exe_rd;
  assign N729 = N728 & fpu1_v_r;
  assign N728 = id_r[19] & N156;
  assign N732 = N731 & fpu1_v_r;
  assign N731 = id_r[18] & N157;
  assign N735 = N734 & fpu1_v_r;
  assign N734 = id_r[17] & N158;
  assign N738 = N737 & mem_ctrl_r[37];
  assign N737 = id_r[19] & id_rs1_equal_mem_rd;
  assign N741 = N740 & mem_ctrl_r[37];
  assign N740 = id_r[18] & id_rs2_equal_mem_rd;
  assign N744 = N743 & mem_ctrl_r[37];
  assign N743 = id_r[17] & id_rs3_equal_mem_rd;
  assign stall_bypass_fp_rs1 = N745 & N754;
  assign N745 = id_r[43] & N651;
  assign N754 = N752 | N753;
  assign N752 = N750 | N751;
  assign N750 = N748 | N749;
  assign N748 = N746 | N747;
  assign N746 = id_rs1_equal_fp_exe_rd & fp_exe_ctrl_r[12];
  assign N747 = N159 & imul_v_lo;
  assign N749 = id_rs1_equal_exe_rd & exe_r[126];
  assign N751 = id_rs1_equal_mem_rd & mem_ctrl_r[38];
  assign N753 = id_rs1_equal_wb_rd & wb_ctrl_r[39];
  assign stall_bypass_int_frs2 = id_r[18] & N763;
  assign N763 = N761 | N762;
  assign N761 = N759 | N760;
  assign N759 = N757 | N758;
  assign N757 = N755 | N756;
  assign N755 = id_rs2_equal_fp_exe_rd & fp_exe_ctrl_r[13];
  assign N756 = N160 & fpu1_v_r;
  assign N758 = N161 & fpu_float_v_lo;
  assign N760 = id_rs2_equal_mem_rd & mem_ctrl_r[37];
  assign N762 = N162 & flw_wb_ctrl_r[5];
  assign N163 = stall_bypass_fp_frs | stall_bypass_fp_rs1;
  assign stall_lr_aq = N765 & N766;
  assign N765 = id_r[27] & N764;
  assign N764 = reserved_r | lsu_reserve_lo;
  assign N766 = ~break_reserve;
  assign stall_fence = id_r[28] & N767;
  assign N767 = N620 | lsu_remote_req_v_lo;
  assign stall_amo_aq = N769 & N773;
  assign N769 = aq_r & N768;
  assign N768 = ~aq_clear;
  assign N773 = N772 | id_r[26];
  assign N772 = N771 | id_r[27];
  assign N771 = N770 | id_r[25];
  assign N770 = id_r[40] | id_r[39];
  assign stall_amo_rl = N774 & N775;
  assign N774 = id_r[25] & id_r[23];
  assign N775 = N620 | lsu_remote_req_v_lo;
  assign local_mem_op_restore = N779 & N780;
  assign N779 = N777 & N778;
  assign N777 = lsu_dmem_v_lo & N776;
  assign N776 = ~exe_r[111];
  assign N778 = ~exe_r[112];
  assign N780 = ~stall_all;
  assign id_remote_req_op = N782 | id_r[1];
  assign N782 = N781 | id_r[25];
  assign N781 = id_r[40] | id_r[39];
  assign memory_op_issued = N785 & N786;
  assign N785 = N783 & N784;
  assign N783 = id_remote_req_op & N684;
  assign N784 = ~stall_id;
  assign N786 = ~stall_all;
  assign N168 = ~reset_i;
  assign stall_remote_req = id_remote_req_op & N171;
  assign stall_remote_credit = id_remote_req_op & N178;
  assign N179 = ~fdiv_fsqrt_ready_lo;
  assign N180 = fp_exe_ctrl_r[11] | fp_exe_ctrl_r[10];
  assign stall_fdiv_busy = N787 & N181;
  assign N787 = id_r[10] | id_r[9];
  assign N182 = ~idiv_ready_lo;
  assign stall_idiv_busy = id_r[31] & N183;
  assign stall_fcsr = N789 & N796;
  assign N789 = id_r[15] & N788;
  assign N788 = N633 | N647;
  assign N796 = N795 | fpu_float_v_lo;
  assign N795 = N794 | fpu1_v_r;
  assign N794 = N793 | fdiv_fsqrt_v_lo;
  assign N793 = N792 | N179;
  assign N792 = N791 | fp_exe_ctrl_r[10];
  assign N791 = N790 | fp_exe_ctrl_r[11];
  assign N790 = fp_exe_ctrl_r[13] | fp_exe_ctrl_r[12];
  assign frs1_forward_v = N797 & float_rf_wen;
  assign N797 = id_r[19] & N184;
  assign frs2_forward_v = N798 & float_rf_wen;
  assign N798 = id_r[18] & N185;
  assign frs3_forward_v = N799 & float_rf_wen;
  assign N799 = id_r[17] & N186;
  assign has_forward_data_rs1[0] = N802 & N651;
  assign N802 = N800 | N801;
  assign N800 = exe_r[126] & id_rs1_equal_exe_rd;
  assign N801 = fp_exe_ctrl_r[12] & id_rs1_equal_fp_exe_rd;
  assign has_forward_data_rs1[1] = N805 & N651;
  assign N805 = N803 | N804;
  assign N803 = mem_ctrl_r[38] & id_rs1_equal_mem_rd;
  assign N804 = imul_v_lo & N187;
  assign has_forward_data_rs1[2] = N806 & N651;
  assign N806 = wb_ctrl_r[39] & id_rs1_equal_wb_rd;
  assign has_forward_data_rs2[0] = N809 & N615;
  assign N809 = N807 | N808;
  assign N807 = exe_r[126] & id_rs2_equal_exe_rd;
  assign N808 = fp_exe_ctrl_r[12] & id_rs2_equal_fp_exe_rd;
  assign has_forward_data_rs2[1] = N812 & N615;
  assign N812 = N810 | N811;
  assign N810 = mem_ctrl_r[38] & id_rs2_equal_mem_rd;
  assign N811 = imul_v_lo & N188;
  assign has_forward_data_rs2[2] = N813 & N615;
  assign N813 = wb_ctrl_r[39] & id_rs2_equal_wb_rd;
  assign aq_set = N817 & N784;
  assign N817 = N815 & N816;
  assign N815 = N814 & N684;
  assign N814 = id_r[25] & id_r[24];
  assign N816 = ~stall_all;
  assign aq_clear = wb_ctrl_r[39] & N189;
  assign fcsr_v_li = N820 & N784;
  assign N820 = N818 & N819;
  assign N818 = id_r[15] & N684;
  assign N819 = ~stall_all;
  assign mcsr_we_li = N823 & N784;
  assign N823 = N821 & N822;
  assign N821 = id_r[15] & N684;
  assign N822 = ~stall_all;
  assign mcsr_instr_executed_li = N827 & mstatus_r_mie_;
  assign N827 = N826 & N784;
  assign N826 = N824 & N825;
  assign N824 = id_r[0] & N684;
  assign N825 = ~stall_all;
  assign mcsr_interrupt_entered_li = interrupt_ready & N828;
  assign N828 = ~stall_all;
  assign mcsr_mret_called_li = exe_r[99] & N829;
  assign N829 = ~stall_all;
  assign N190 = ~stall_all;
  assign N191 = stall_all;
  assign N192 = N830 | exe_r[99];
  assign N830 = exe_r[0] & mstatus_r_mie_;
  assign N193 = flush | stall_id;
  assign N194 = id_r[20] | N193;
  assign N195 = ~N194;
  assign N196 = ~id_r[15];
  assign N197 = ~fcsr_data_v_lo;
  assign N487 = ~N193;
  assign N488 = id_r[20] & N487;
  assign idiv_v_li = exe_r[116] & N831;
  assign N831 = ~stall_all;
  assign int_sb_score = N832 & N834;
  assign N832 = ~stall_all;
  assign N834 = N833 | int_remote_load_in_exe;
  assign N833 = exe_r[116] | exe_r[110];
  assign N489 = ~fp_exe_ctrl_r[12];
  assign remote_req_v_o = lsu_remote_req_v_lo & N835;
  assign N835 = ~stall_all;
  assign N490 = ~N611;
  assign N491 = N836 | N837;
  assign N836 = flush | stall_id;
  assign N837 = ~id_r[20];
  assign N492 = stall_all;
  assign N493 = N491 | N492;
  assign N494 = ~N493;
  assign N495 = N493;
  assign N496 = ~N492;
  assign N497 = N491 & N496;
  assign fdiv_fsqrt_v_li = fdiv_fsqrt_in_fp_exe & N838;
  assign N838 = ~stall_all;
  assign float_sb_score = N839 & N840;
  assign N839 = ~stall_all;
  assign N840 = fdiv_fsqrt_in_fp_exe | float_remote_load_in_exe;
  assign N498 = ~fdiv_fsqrt_in_fp_exe;
  assign N499 = exe_r[116] | N842;
  assign N842 = lsu_remote_req_v_lo & N841;
  assign N841 = ~exe_r[1];
  assign N500 = stall_all;
  assign N501 = N499 | N500;
  assign N502 = fp_exe_ctrl_r[12] | N501;
  assign N503 = ~N502;
  assign N504 = ~N500;
  assign N505 = N499 & N504;
  assign N506 = ~N499;
  assign N507 = N504 & N506;
  assign N508 = fp_exe_ctrl_r[12] & N507;
  assign N509 = stall_all;
  assign N510 = lsu_dmem_v_lo | N509;
  assign N511 = ~N510;
  assign N512 = ~N509;
  assign N513 = lsu_dmem_v_lo & N512;
  assign make_reserve = lsu_reserve_lo & N843;
  assign N843 = ~stall_all;
  assign break_reserve = N845 & dmem_w_li;
  assign N845 = N844 & dmem_v_li;
  assign N844 = reserved_r & N514;
  assign stall_ifetch_wait = mem_ctrl_r[0] & N132;
  assign N515 = mem_ctrl_r[33] | imul_v_lo;
  assign N516 = ~N515;
  assign N517 = ~imul_v_lo;
  assign N518 = mem_ctrl_r[33] & N517;
  assign mem_result_valid = N846 | mem_ctrl_r[37];
  assign N846 = imul_v_lo | mem_ctrl_r[38];
  assign N519 = mem_ctrl_r[0] & ifetch_v_i;
  assign N520 = N519 | int_remote_load_resp_force_i;
  assign N521 = imul_v_lo | N520;
  assign N522 = mem_ctrl_r[38] | N521;
  assign N523 = int_remote_load_resp_v_i | N522;
  assign N524 = idiv_v_lo | N523;
  assign N525 = ~N524;
  assign N526 = mem_result_valid | mem_ctrl_r[0];
  assign N527 = ~mem_ctrl_r[33];
  assign N560 = ~wb_ctrl_n[33];
  assign N561 = N560;
  assign N562 = ~int_remote_load_resp_force_i;
  assign N563 = ~N523;
  assign wb_ctrl_n[33] = N519 & N562;
  assign N564 = ~N519;
  assign N565 = N562 & N564;
  assign N566 = imul_v_lo & N565;
  assign N567 = N565 & N517;
  assign N568 = mem_ctrl_r[38] & N567;
  assign N569 = ~mem_ctrl_r[38];
  assign N570 = N567 & N569;
  assign N571 = int_remote_load_resp_v_i & N570;
  assign N572 = ~int_remote_load_resp_v_i;
  assign N573 = N570 & N572;
  assign N574 = idiv_v_lo & N573;
  assign int_sb_clear = wb_ctrl_r[39] & wb_ctrl_r[0];
  assign N575 = ~stall_all;
  assign N576 = stall_all;
  assign N577 = flw_wb_ctrl_r[5] | float_remote_load_resp_force_i;
  assign N578 = fpu_float_v_lo | N577;
  assign N579 = fdiv_fsqrt_v_lo | N578;
  assign N580 = float_remote_load_resp_v_i | N579;
  assign N581 = ~N580;
  assign N582 = flw_wb_ctrl_r[5] | fpu_float_v_lo;
  assign N583 = ~float_remote_load_resp_force_i;
  assign N584 = ~N593;
  assign N585 = N584;
  assign N586 = ~N579;
  assign N587 = flw_wb_ctrl_r[5] & N583;
  assign N588 = ~flw_wb_ctrl_r[5];
  assign N589 = N583 & N588;
  assign N590 = fpu_float_v_lo & N589;
  assign N591 = ~fpu_float_v_lo;
  assign N592 = N589 & N591;
  assign N593 = fdiv_fsqrt_v_lo & N592;
  assign N594 = ~fdiv_fsqrt_v_lo;
  assign N595 = N592 & N594;
  assign N596 = float_remote_load_resp_v_i & N595;
  assign stall_fpu2_li = 1'b0 | stall_remote_flw_wb;

  always @(posedge clk_i) begin
    if(reset_i) begin
      aq_rd_r_4_sv2v_reg <= 1'b0;
      aq_rd_r_3_sv2v_reg <= 1'b0;
      aq_rd_r_2_sv2v_reg <= 1'b0;
      aq_rd_r_1_sv2v_reg <= 1'b0;
      aq_rd_r_0_sv2v_reg <= 1'b0;
    end else if(N47) begin
      aq_rd_r_4_sv2v_reg <= id_r[55];
      aq_rd_r_3_sv2v_reg <= id_r[54];
      aq_rd_r_2_sv2v_reg <= id_r[53];
      aq_rd_r_1_sv2v_reg <= id_r[52];
      aq_rd_r_0_sv2v_reg <= id_r[51];
    end 
    if(reset_i) begin
      aq_r_sv2v_reg <= 1'b0;
    end else if(N46) begin
      aq_r_sv2v_reg <= aq_set;
    end 
    if(reset_i) begin
      reserved_addr_r_9_sv2v_reg <= 1'b0;
      reserved_addr_r_8_sv2v_reg <= 1'b0;
      reserved_addr_r_7_sv2v_reg <= 1'b0;
      reserved_addr_r_6_sv2v_reg <= 1'b0;
      reserved_addr_r_5_sv2v_reg <= 1'b0;
      reserved_addr_r_4_sv2v_reg <= 1'b0;
      reserved_addr_r_3_sv2v_reg <= 1'b0;
      reserved_addr_r_2_sv2v_reg <= 1'b0;
      reserved_addr_r_1_sv2v_reg <= 1'b0;
      reserved_addr_r_0_sv2v_reg <= 1'b0;
    end else if(N73) begin
      reserved_addr_r_9_sv2v_reg <= dmem_addr_li[9];
      reserved_addr_r_8_sv2v_reg <= dmem_addr_li[8];
      reserved_addr_r_7_sv2v_reg <= dmem_addr_li[7];
      reserved_addr_r_6_sv2v_reg <= dmem_addr_li[6];
      reserved_addr_r_5_sv2v_reg <= dmem_addr_li[5];
      reserved_addr_r_4_sv2v_reg <= dmem_addr_li[4];
      reserved_addr_r_3_sv2v_reg <= dmem_addr_li[3];
      reserved_addr_r_2_sv2v_reg <= dmem_addr_li[2];
      reserved_addr_r_1_sv2v_reg <= dmem_addr_li[1];
      reserved_addr_r_0_sv2v_reg <= dmem_addr_li[0];
    end 
    if(reset_i) begin
      reserved_r_sv2v_reg <= 1'b0;
    end else if(N72) begin
      reserved_r_sv2v_reg <= make_reserve;
    end 
    if(reset_i) begin
      remote_req_counter_r_1_sv2v_reg <= 1'b1;
      remote_req_counter_r_0_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      remote_req_counter_r_1_sv2v_reg <= N170;
      remote_req_counter_r_0_sv2v_reg <= N169;
    end 
  end


endmodule



module bsg_manycore_proc_vanilla_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_data_width_p32_addr_width_p28_icache_tag_width_p12_icache_entries_p1024_dmem_size_p1024_num_vcache_rows_p1_vcache_size_pinv_vcache_sets_pinv_num_tiles_x_p16_num_tiles_y_p8_rev_fifo_els_p2_fwd_fifo_els_p3_debug_p0
(
  clk_i,
  reset_i,
  link_sif_i,
  link_sif_o,
  my_x_i,
  my_y_i,
  pod_x_i,
  pod_y_i
);

  input [153:0] link_sif_i;
  output [153:0] link_sif_o;
  input [3:0] my_x_i;
  input [2:0] my_y_i;
  input [2:0] pod_x_i;
  input [3:0] pod_y_i;
  input clk_i;
  input reset_i;
  wire [153:0] link_sif_o;
  wire in_v_lo,in_we_lo,in_yumi_li,returning_data_v_li,out_v_li,out_credit_or_ready_lo,
  returned_v_r_lo,returned_fifo_full_lo,returned_yumi_li,remote_dmem_v_lo,
  remote_dmem_w_lo,remote_dmem_yumi_li,icache_v_lo,icache_yumi_li,freeze,
  remote_interrupt_set_lo,remote_interrupt_clear_lo,remote_interrupt_pending_bit_li,remote_req_v,
  remote_req_credit,ifetch_v_lo,float_remote_load_resp_v_lo,
  float_remote_load_resp_force_lo,float_remote_load_resp_yumi_li,int_remote_load_resp_v_lo,
  int_remote_load_resp_force_lo,int_remote_load_resp_yumi_li,invalid_eva_access_lo,sv2v_dc_1,
  sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5;
  wire [27:0] in_addr_lo;
  wire [31:0] in_data_lo,returning_data_li,returned_data_r_lo,remote_dmem_data_lo,
  remote_dmem_data_li,icache_instr_lo,ifetch_instr_lo,float_remote_load_resp_data_lo,
  int_remote_load_resp_data_lo;
  wire [3:0] in_mask_lo,remote_dmem_mask_lo,tgo_x,cfg_pod_y_lo;
  wire [6:0] in_load_info_lo,src_x_cord_debug_lo,src_y_cord_debug_lo;
  wire [96:0] out_packet_li;
  wire [4:0] returned_reg_id_r_lo,float_remote_load_resp_rd_lo,int_remote_load_resp_rd_lo;
  wire [1:0] returned_pkt_type_r_lo;
  wire [5:0] out_credits_used_lo;
  wire [9:0] remote_dmem_addr_lo;
  wire [21:0] icache_pc_lo,pc_init_val;
  wire [2:0] tgo_y,cfg_pod_x_lo;
  wire [83:0] remote_req;

  bsg_manycore_endpoint_standard_x_cord_width_p7_y_cord_width_p7_fifo_els_p4_data_width_p32_addr_width_p28_credit_counter_width_p6_rev_fifo_els_p2_use_credits_for_local_fifo_p1
  endp
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_sif_i(link_sif_i),
    .link_sif_o(link_sif_o),
    .in_v_o(in_v_lo),
    .in_data_o(in_data_lo),
    .in_mask_o(in_mask_lo),
    .in_addr_o(in_addr_lo),
    .in_we_o(in_we_lo),
    .in_load_info_o(in_load_info_lo),
    .in_src_x_cord_o(src_x_cord_debug_lo),
    .in_src_y_cord_o(src_y_cord_debug_lo),
    .in_yumi_i(in_yumi_li),
    .returning_data_i(returning_data_li),
    .returning_v_i(returning_data_v_li),
    .out_v_i(out_v_li),
    .out_packet_i(out_packet_li),
    .out_credit_or_ready_o(out_credit_or_ready_lo),
    .returned_data_r_o(returned_data_r_lo),
    .returned_reg_id_r_o(returned_reg_id_r_lo),
    .returned_v_r_o(returned_v_r_lo),
    .returned_pkt_type_r_o(returned_pkt_type_r_lo),
    .returned_yumi_i(returned_yumi_li),
    .returned_fifo_full_o(returned_fifo_full_lo),
    .returned_credit_reg_id_r_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5 }),
    .out_credits_used_o(out_credits_used_lo),
    .global_x_i({ pod_x_i, my_x_i }),
    .global_y_i({ pod_y_i, my_y_i })
  );


  network_rx_data_width_p32_addr_width_p28_dmem_size_p1024_icache_tag_width_p12_icache_entries_p1024_x_cord_width_p7_y_cord_width_p7_x_subcord_width_p4_y_subcord_width_p3
  rx
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(in_v_lo),
    .w_i(in_we_lo),
    .addr_i(in_addr_lo),
    .data_i(in_data_lo),
    .mask_i(in_mask_lo),
    .load_info_i(in_load_info_lo),
    .yumi_o(in_yumi_li),
    .src_x_cord_debug_i(src_x_cord_debug_lo),
    .src_y_cord_debug_i(src_y_cord_debug_lo),
    .returning_data_o(returning_data_li),
    .returning_data_v_o(returning_data_v_li),
    .remote_dmem_v_o(remote_dmem_v_lo),
    .remote_dmem_w_o(remote_dmem_w_lo),
    .remote_dmem_addr_o(remote_dmem_addr_lo),
    .remote_dmem_mask_o(remote_dmem_mask_lo),
    .remote_dmem_data_o(remote_dmem_data_lo),
    .remote_dmem_data_i(remote_dmem_data_li),
    .remote_dmem_yumi_i(remote_dmem_yumi_li),
    .icache_v_o(icache_v_lo),
    .icache_pc_o(icache_pc_lo),
    .icache_instr_o(icache_instr_lo),
    .icache_yumi_i(icache_yumi_li),
    .freeze_o(freeze),
    .tgo_x_o(tgo_x),
    .tgo_y_o(tgo_y),
    .pc_init_val_o(pc_init_val),
    .remote_interrupt_set_o(remote_interrupt_set_lo),
    .remote_interrupt_clear_o(remote_interrupt_clear_lo),
    .remote_interrupt_pending_bit_i(remote_interrupt_pending_bit_li),
    .global_x_i({ pod_x_i, my_x_i }),
    .global_y_i({ pod_y_i, my_y_i })
  );


  network_tx_data_width_p32_addr_width_p28_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_num_vcache_rows_p1_vcache_size_pinv_vcache_sets_pinv_num_tiles_x_p16_num_tiles_y_p8_icache_entries_p1024_icache_tag_width_p12
  tx
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .out_packet_o(out_packet_li),
    .out_v_o(out_v_li),
    .out_credit_or_ready_i(out_credit_or_ready_lo),
    .returned_v_i(returned_v_r_lo),
    .returned_data_i(returned_data_r_lo),
    .returned_reg_id_i(returned_reg_id_r_lo),
    .returned_pkt_type_i(returned_pkt_type_r_lo),
    .returned_fifo_full_i(returned_fifo_full_lo),
    .returned_yumi_o(returned_yumi_li),
    .tgo_x_i(tgo_x),
    .tgo_y_i(tgo_y),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .pod_x_i(pod_x_i),
    .pod_y_i(pod_y_i),
    .cfg_pod_x_i(cfg_pod_x_lo),
    .cfg_pod_y_i(cfg_pod_y_lo),
    .remote_req_i(remote_req),
    .remote_req_v_i(remote_req_v),
    .remote_req_credit_o(remote_req_credit),
    .ifetch_v_o(ifetch_v_lo),
    .ifetch_instr_o(ifetch_instr_lo),
    .float_remote_load_resp_rd_o(float_remote_load_resp_rd_lo),
    .float_remote_load_resp_data_o(float_remote_load_resp_data_lo),
    .float_remote_load_resp_v_o(float_remote_load_resp_v_lo),
    .float_remote_load_resp_force_o(float_remote_load_resp_force_lo),
    .float_remote_load_resp_yumi_i(float_remote_load_resp_yumi_li),
    .int_remote_load_resp_rd_o(int_remote_load_resp_rd_lo),
    .int_remote_load_resp_data_o(int_remote_load_resp_data_lo),
    .int_remote_load_resp_v_o(int_remote_load_resp_v_lo),
    .int_remote_load_resp_force_o(int_remote_load_resp_force_lo),
    .int_remote_load_resp_yumi_i(int_remote_load_resp_yumi_li),
    .invalid_eva_access_o(invalid_eva_access_lo)
  );


  vanilla_core_data_width_p32_dmem_size_p1024_icache_entries_p1024_icache_tag_width_p12_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_credit_counter_width_p6_fwd_fifo_els_p3
  vcore
  (
    .clk_i(clk_i),
    .reset_i(freeze),
    .pc_init_val_i(pc_init_val),
    .remote_req_o(remote_req),
    .remote_req_v_o(remote_req_v),
    .remote_req_credit_i(remote_req_credit),
    .icache_v_i(icache_v_lo),
    .icache_pc_i(icache_pc_lo),
    .icache_instr_i(icache_instr_lo),
    .icache_yumi_o(icache_yumi_li),
    .ifetch_v_i(ifetch_v_lo),
    .ifetch_instr_i(ifetch_instr_lo),
    .remote_dmem_v_i(remote_dmem_v_lo),
    .remote_dmem_w_i(remote_dmem_w_lo),
    .remote_dmem_addr_i(remote_dmem_addr_lo),
    .remote_dmem_mask_i(remote_dmem_mask_lo),
    .remote_dmem_data_i(remote_dmem_data_lo),
    .remote_dmem_data_o(remote_dmem_data_li),
    .remote_dmem_yumi_o(remote_dmem_yumi_li),
    .float_remote_load_resp_rd_i(float_remote_load_resp_rd_lo),
    .float_remote_load_resp_data_i(float_remote_load_resp_data_lo),
    .float_remote_load_resp_v_i(float_remote_load_resp_v_lo),
    .float_remote_load_resp_force_i(float_remote_load_resp_force_lo),
    .float_remote_load_resp_yumi_o(float_remote_load_resp_yumi_li),
    .int_remote_load_resp_rd_i(int_remote_load_resp_rd_lo),
    .int_remote_load_resp_data_i(int_remote_load_resp_data_lo),
    .int_remote_load_resp_v_i(int_remote_load_resp_v_lo),
    .int_remote_load_resp_force_i(int_remote_load_resp_force_lo),
    .int_remote_load_resp_yumi_o(int_remote_load_resp_yumi_li),
    .invalid_eva_access_i(invalid_eva_access_lo),
    .remote_interrupt_set_i(remote_interrupt_set_lo),
    .remote_interrupt_clear_i(remote_interrupt_clear_lo),
    .remote_interrupt_pending_bit_o(remote_interrupt_pending_bit_li),
    .out_credits_used_i(out_credits_used_lo),
    .cfg_pod_x_o(cfg_pod_x_lo),
    .cfg_pod_y_o(cfg_pod_y_lo),
    .global_x_i({ pod_x_i, my_x_i }),
    .global_y_i({ pod_y_i, my_y_i })
  );


endmodule



module bsg_manycore_hetero_socket_x_cord_width_p7_y_cord_width_p7_data_width_p32_addr_width_p28_dmem_size_p1024_icache_entries_p1024_icache_tag_width_p12_num_vcache_rows_p1_vcache_size_pinv_debug_p0_hetero_type_p0_pod_x_cord_width_p3_pod_y_cord_width_p4_num_tiles_x_p16_num_tiles_y_p8_vcache_sets_pinv_fwd_fifo_els_p3_rev_fifo_els_p2
(
  clk_i,
  reset_i,
  link_sif_i,
  link_sif_o,
  my_x_i,
  my_y_i,
  pod_x_i,
  pod_y_i
);

  input [153:0] link_sif_i;
  output [153:0] link_sif_o;
  input [3:0] my_x_i;
  input [2:0] my_y_i;
  input [2:0] pod_x_i;
  input [3:0] pod_y_i;
  input clk_i;
  input reset_i;
  wire [153:0] link_sif_o;

  bsg_manycore_proc_vanilla_x_cord_width_p7_y_cord_width_p7_pod_x_cord_width_p3_pod_y_cord_width_p4_data_width_p32_addr_width_p28_icache_tag_width_p12_icache_entries_p1024_dmem_size_p1024_num_vcache_rows_p1_vcache_size_pinv_vcache_sets_pinv_num_tiles_x_p16_num_tiles_y_p8_rev_fifo_els_p2_fwd_fifo_els_p3_debug_p0
  \h.z 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_sif_i(link_sif_i),
    .link_sif_o(link_sif_o),
    .my_x_i(my_x_i),
    .my_y_i(my_y_i),
    .pod_x_i(pod_x_i),
    .pod_y_i(pod_y_i)
  );


endmodule



module bsg_manycore_withfakeram
(
  clk_i,
  reset_i,
  reset_o,
  link_i,
  link_o,
  global_x_i,
  global_y_i,
  global_x_o,
  global_y_o
);

  input [615:0] link_i;
  output [615:0] link_o;
  input [6:0] global_x_i;
  input [6:0] global_y_i;
  output [6:0] global_x_o;
  output [6:0] global_y_o;
  input clk_i;
  input reset_i;
  output reset_o;
  wire [615:0] link_o;
  wire [6:0] global_x_o,global_y_o;
  wire reset_o,reset_r;
  wire [3:0] pod_y_r;
  wire [2:0] my_y_r;
  wire [153:0] proc_link_sif_li,proc_link_sif_lo;

  bsg_dff_width_p1
  dff_reset
  (
    .clk_i(clk_i),
    .data_i(reset_i),
    .data_o(reset_r)
  );


  bsg_dff_width_p7
  dff_x
  (
    .clk_i(clk_i),
    .data_i(global_x_i),
    .data_o(global_x_o)
  );


  bsg_dff_width_p7
  dff_y
  (
    .clk_i(clk_i),
    .data_i(global_y_i),
    .data_o({ pod_y_r, my_y_r })
  );


  bsg_manycore_mesh_node_7_7_32_28_2_0_0_01_00_0
  rtr
  (
    .clk_i(clk_i),
    .reset_i(reset_r),
    .links_sif_i(link_i),
    .links_sif_o(link_o),
    .proc_link_sif_i(proc_link_sif_li),
    .proc_link_sif_o(proc_link_sif_lo),
    .global_x_i(global_x_o),
    .global_y_i({ pod_y_r, my_y_r })
  );


  bsg_manycore_hetero_socket_x_cord_width_p7_y_cord_width_p7_data_width_p32_addr_width_p28_dmem_size_p1024_icache_entries_p1024_icache_tag_width_p12_num_vcache_rows_p1_vcache_size_pinv_debug_p0_hetero_type_p0_pod_x_cord_width_p3_pod_y_cord_width_p4_num_tiles_x_p16_num_tiles_y_p8_vcache_sets_pinv_fwd_fifo_els_p3_rev_fifo_els_p2
  proc
  (
    .clk_i(clk_i),
    .reset_i(reset_r),
    .link_sif_i(proc_link_sif_lo),
    .link_sif_o(proc_link_sif_li),
    .my_x_i(global_x_o[3:0]),
    .my_y_i(my_y_r),
    .pod_x_i(global_x_o[6:4]),
    .pod_y_i(pod_y_r)
  );

  assign global_y_o = { pod_y_r, my_y_r } + 1'b1;

endmodule

