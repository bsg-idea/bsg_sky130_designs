VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_64x96
  FOREIGN fakeram130_64x96 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1800.000 BY 800.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.550 0.900 18.450 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 19.350 0.900 20.250 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.150 0.900 22.050 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.950 0.900 23.850 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.750 0.900 25.650 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.550 0.900 27.450 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.350 0.900 29.250 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 30.150 0.900 31.050 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.950 0.900 32.850 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.750 0.900 34.650 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.550 0.900 36.450 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.350 0.900 38.250 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.150 0.900 40.050 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.950 0.900 41.850 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.750 0.900 43.650 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.550 0.900 45.450 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 46.350 0.900 47.250 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 48.150 0.900 49.050 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 49.950 0.900 50.850 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 51.750 0.900 52.650 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 53.550 0.900 54.450 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.350 0.900 56.250 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 57.150 0.900 58.050 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 58.950 0.900 59.850 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 60.750 0.900 61.650 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.550 0.900 63.450 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.350 0.900 65.250 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.150 0.900 67.050 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.950 0.900 68.850 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.750 0.900 70.650 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.550 0.900 72.450 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.350 0.900 74.250 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 75.150 0.900 76.050 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.950 0.900 77.850 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.750 0.900 79.650 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.550 0.900 81.450 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.350 0.900 83.250 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.150 0.900 85.050 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.950 0.900 86.850 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 87.750 0.900 88.650 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.550 0.900 90.450 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 91.350 0.900 92.250 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.150 0.900 94.050 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.950 0.900 95.850 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.750 0.900 97.650 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 98.550 0.900 99.450 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.350 0.900 101.250 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.150 0.900 103.050 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.950 0.900 104.850 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.750 0.900 106.650 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.550 0.900 108.450 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 109.350 0.900 110.250 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.150 0.900 112.050 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.950 0.900 113.850 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 114.750 0.900 115.650 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.550 0.900 117.450 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.350 0.900 119.250 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.150 0.900 121.050 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 121.950 0.900 122.850 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.750 0.900 124.650 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 125.550 0.900 126.450 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.350 0.900 128.250 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 129.150 0.900 130.050 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.950 0.900 131.850 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 132.750 0.900 133.650 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.550 0.900 135.450 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.350 0.900 137.250 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 138.150 0.900 139.050 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.950 0.900 140.850 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.750 0.900 142.650 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.550 0.900 144.450 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.350 0.900 146.250 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 147.150 0.900 148.050 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.950 0.900 149.850 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.750 0.900 151.650 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.550 0.900 153.450 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.350 0.900 155.250 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.150 0.900 157.050 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.950 0.900 158.850 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 159.750 0.900 160.650 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.550 0.900 162.450 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.350 0.900 164.250 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.150 0.900 166.050 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.950 0.900 167.850 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.750 0.900 169.650 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 170.550 0.900 171.450 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 172.350 0.900 173.250 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 174.150 0.900 175.050 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 175.950 0.900 176.850 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 177.750 0.900 178.650 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 179.550 0.900 180.450 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 181.350 0.900 182.250 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 183.150 0.900 184.050 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 184.950 0.900 185.850 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 186.750 0.900 187.650 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 188.550 0.900 189.450 ;
    END
  END w_mask_in[95]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 244.350 0.900 245.250 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 246.150 0.900 247.050 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 247.950 0.900 248.850 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 249.750 0.900 250.650 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 251.550 0.900 252.450 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 253.350 0.900 254.250 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 255.150 0.900 256.050 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 256.950 0.900 257.850 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 258.750 0.900 259.650 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 260.550 0.900 261.450 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 262.350 0.900 263.250 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 264.150 0.900 265.050 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 265.950 0.900 266.850 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 267.750 0.900 268.650 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 269.550 0.900 270.450 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 271.350 0.900 272.250 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 273.150 0.900 274.050 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 274.950 0.900 275.850 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 276.750 0.900 277.650 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 278.550 0.900 279.450 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 280.350 0.900 281.250 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 282.150 0.900 283.050 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 283.950 0.900 284.850 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 285.750 0.900 286.650 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 287.550 0.900 288.450 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 289.350 0.900 290.250 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 291.150 0.900 292.050 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 292.950 0.900 293.850 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 294.750 0.900 295.650 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 296.550 0.900 297.450 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 298.350 0.900 299.250 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 300.150 0.900 301.050 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 301.950 0.900 302.850 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 303.750 0.900 304.650 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 305.550 0.900 306.450 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 307.350 0.900 308.250 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 309.150 0.900 310.050 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 310.950 0.900 311.850 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 312.750 0.900 313.650 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 314.550 0.900 315.450 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 316.350 0.900 317.250 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 318.150 0.900 319.050 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 319.950 0.900 320.850 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 321.750 0.900 322.650 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 323.550 0.900 324.450 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 325.350 0.900 326.250 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.150 0.900 328.050 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 328.950 0.900 329.850 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.750 0.900 331.650 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 332.550 0.900 333.450 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 334.350 0.900 335.250 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 336.150 0.900 337.050 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.950 0.900 338.850 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 339.750 0.900 340.650 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 341.550 0.900 342.450 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 343.350 0.900 344.250 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 345.150 0.900 346.050 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 346.950 0.900 347.850 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 348.750 0.900 349.650 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 350.550 0.900 351.450 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 352.350 0.900 353.250 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 354.150 0.900 355.050 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 355.950 0.900 356.850 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 357.750 0.900 358.650 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 359.550 0.900 360.450 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 361.350 0.900 362.250 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 363.150 0.900 364.050 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 364.950 0.900 365.850 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 366.750 0.900 367.650 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 368.550 0.900 369.450 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 370.350 0.900 371.250 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 372.150 0.900 373.050 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 373.950 0.900 374.850 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 375.750 0.900 376.650 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 377.550 0.900 378.450 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 379.350 0.900 380.250 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 381.150 0.900 382.050 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 382.950 0.900 383.850 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 384.750 0.900 385.650 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 386.550 0.900 387.450 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 388.350 0.900 389.250 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 390.150 0.900 391.050 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 391.950 0.900 392.850 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 393.750 0.900 394.650 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 395.550 0.900 396.450 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 397.350 0.900 398.250 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.150 0.900 400.050 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 400.950 0.900 401.850 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 402.750 0.900 403.650 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 404.550 0.900 405.450 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 406.350 0.900 407.250 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 408.150 0.900 409.050 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.950 0.900 410.850 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 411.750 0.900 412.650 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 413.550 0.900 414.450 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 415.350 0.900 416.250 ;
    END
  END rd_out[95]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 471.150 0.900 472.050 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 472.950 0.900 473.850 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 474.750 0.900 475.650 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 476.550 0.900 477.450 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 478.350 0.900 479.250 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 480.150 0.900 481.050 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 481.950 0.900 482.850 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 483.750 0.900 484.650 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.550 0.900 486.450 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 487.350 0.900 488.250 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 489.150 0.900 490.050 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 490.950 0.900 491.850 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 492.750 0.900 493.650 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 494.550 0.900 495.450 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 496.350 0.900 497.250 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 498.150 0.900 499.050 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 499.950 0.900 500.850 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.750 0.900 502.650 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 503.550 0.900 504.450 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 505.350 0.900 506.250 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 507.150 0.900 508.050 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 508.950 0.900 509.850 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 510.750 0.900 511.650 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 512.550 0.900 513.450 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 514.350 0.900 515.250 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 516.150 0.900 517.050 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 517.950 0.900 518.850 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 519.750 0.900 520.650 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 521.550 0.900 522.450 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 523.350 0.900 524.250 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 525.150 0.900 526.050 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.950 0.900 527.850 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 528.750 0.900 529.650 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 530.550 0.900 531.450 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 532.350 0.900 533.250 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 534.150 0.900 535.050 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.950 0.900 536.850 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 537.750 0.900 538.650 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 539.550 0.900 540.450 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 541.350 0.900 542.250 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.150 0.900 544.050 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 544.950 0.900 545.850 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 546.750 0.900 547.650 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 548.550 0.900 549.450 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 550.350 0.900 551.250 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 552.150 0.900 553.050 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 553.950 0.900 554.850 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 555.750 0.900 556.650 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 557.550 0.900 558.450 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 559.350 0.900 560.250 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 561.150 0.900 562.050 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 562.950 0.900 563.850 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 564.750 0.900 565.650 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 566.550 0.900 567.450 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 568.350 0.900 569.250 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 570.150 0.900 571.050 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 571.950 0.900 572.850 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 573.750 0.900 574.650 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 575.550 0.900 576.450 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 577.350 0.900 578.250 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 579.150 0.900 580.050 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 580.950 0.900 581.850 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 582.750 0.900 583.650 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 584.550 0.900 585.450 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 586.350 0.900 587.250 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 588.150 0.900 589.050 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 589.950 0.900 590.850 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 591.750 0.900 592.650 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 593.550 0.900 594.450 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 595.350 0.900 596.250 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 597.150 0.900 598.050 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 598.950 0.900 599.850 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 600.750 0.900 601.650 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 602.550 0.900 603.450 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 604.350 0.900 605.250 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 606.150 0.900 607.050 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 607.950 0.900 608.850 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 609.750 0.900 610.650 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 611.550 0.900 612.450 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 613.350 0.900 614.250 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 615.150 0.900 616.050 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 616.950 0.900 617.850 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 618.750 0.900 619.650 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 620.550 0.900 621.450 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 622.350 0.900 623.250 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 624.150 0.900 625.050 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 625.950 0.900 626.850 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 627.750 0.900 628.650 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 629.550 0.900 630.450 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 631.350 0.900 632.250 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 633.150 0.900 634.050 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 634.950 0.900 635.850 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 636.750 0.900 637.650 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 638.550 0.900 639.450 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 640.350 0.900 641.250 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 642.150 0.900 643.050 ;
    END
  END wd_in[95]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 697.950 0.900 698.850 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 699.750 0.900 700.650 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 701.550 0.900 702.450 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 703.350 0.900 704.250 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 705.150 0.900 706.050 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 706.950 0.900 707.850 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 762.750 0.900 763.650 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 764.550 0.900 765.450 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 766.350 0.900 767.250 ;
    END
  END clk
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 16.200 18.000 19.800 782.000 ;
      RECT 45.000 18.000 48.600 782.000 ;
      RECT 73.800 18.000 77.400 782.000 ;
      RECT 102.600 18.000 106.200 782.000 ;
      RECT 131.400 18.000 135.000 782.000 ;
      RECT 160.200 18.000 163.800 782.000 ;
      RECT 189.000 18.000 192.600 782.000 ;
      RECT 217.800 18.000 221.400 782.000 ;
      RECT 246.600 18.000 250.200 782.000 ;
      RECT 275.400 18.000 279.000 782.000 ;
      RECT 304.200 18.000 307.800 782.000 ;
      RECT 333.000 18.000 336.600 782.000 ;
      RECT 361.800 18.000 365.400 782.000 ;
      RECT 390.600 18.000 394.200 782.000 ;
      RECT 419.400 18.000 423.000 782.000 ;
      RECT 448.200 18.000 451.800 782.000 ;
      RECT 477.000 18.000 480.600 782.000 ;
      RECT 505.800 18.000 509.400 782.000 ;
      RECT 534.600 18.000 538.200 782.000 ;
      RECT 563.400 18.000 567.000 782.000 ;
      RECT 592.200 18.000 595.800 782.000 ;
      RECT 621.000 18.000 624.600 782.000 ;
      RECT 649.800 18.000 653.400 782.000 ;
      RECT 678.600 18.000 682.200 782.000 ;
      RECT 707.400 18.000 711.000 782.000 ;
      RECT 736.200 18.000 739.800 782.000 ;
      RECT 765.000 18.000 768.600 782.000 ;
      RECT 793.800 18.000 797.400 782.000 ;
      RECT 822.600 18.000 826.200 782.000 ;
      RECT 851.400 18.000 855.000 782.000 ;
      RECT 880.200 18.000 883.800 782.000 ;
      RECT 909.000 18.000 912.600 782.000 ;
      RECT 937.800 18.000 941.400 782.000 ;
      RECT 966.600 18.000 970.200 782.000 ;
      RECT 995.400 18.000 999.000 782.000 ;
      RECT 1024.200 18.000 1027.800 782.000 ;
      RECT 1053.000 18.000 1056.600 782.000 ;
      RECT 1081.800 18.000 1085.400 782.000 ;
      RECT 1110.600 18.000 1114.200 782.000 ;
      RECT 1139.400 18.000 1143.000 782.000 ;
      RECT 1168.200 18.000 1171.800 782.000 ;
      RECT 1197.000 18.000 1200.600 782.000 ;
      RECT 1225.800 18.000 1229.400 782.000 ;
      RECT 1254.600 18.000 1258.200 782.000 ;
      RECT 1283.400 18.000 1287.000 782.000 ;
      RECT 1312.200 18.000 1315.800 782.000 ;
      RECT 1341.000 18.000 1344.600 782.000 ;
      RECT 1369.800 18.000 1373.400 782.000 ;
      RECT 1398.600 18.000 1402.200 782.000 ;
      RECT 1427.400 18.000 1431.000 782.000 ;
      RECT 1456.200 18.000 1459.800 782.000 ;
      RECT 1485.000 18.000 1488.600 782.000 ;
      RECT 1513.800 18.000 1517.400 782.000 ;
      RECT 1542.600 18.000 1546.200 782.000 ;
      RECT 1571.400 18.000 1575.000 782.000 ;
      RECT 1600.200 18.000 1603.800 782.000 ;
      RECT 1629.000 18.000 1632.600 782.000 ;
      RECT 1657.800 18.000 1661.400 782.000 ;
      RECT 1686.600 18.000 1690.200 782.000 ;
      RECT 1715.400 18.000 1719.000 782.000 ;
      RECT 1744.200 18.000 1747.800 782.000 ;
      RECT 1773.000 18.000 1776.600 782.000 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 30.600 18.000 34.200 782.000 ;
      RECT 59.400 18.000 63.000 782.000 ;
      RECT 88.200 18.000 91.800 782.000 ;
      RECT 117.000 18.000 120.600 782.000 ;
      RECT 145.800 18.000 149.400 782.000 ;
      RECT 174.600 18.000 178.200 782.000 ;
      RECT 203.400 18.000 207.000 782.000 ;
      RECT 232.200 18.000 235.800 782.000 ;
      RECT 261.000 18.000 264.600 782.000 ;
      RECT 289.800 18.000 293.400 782.000 ;
      RECT 318.600 18.000 322.200 782.000 ;
      RECT 347.400 18.000 351.000 782.000 ;
      RECT 376.200 18.000 379.800 782.000 ;
      RECT 405.000 18.000 408.600 782.000 ;
      RECT 433.800 18.000 437.400 782.000 ;
      RECT 462.600 18.000 466.200 782.000 ;
      RECT 491.400 18.000 495.000 782.000 ;
      RECT 520.200 18.000 523.800 782.000 ;
      RECT 549.000 18.000 552.600 782.000 ;
      RECT 577.800 18.000 581.400 782.000 ;
      RECT 606.600 18.000 610.200 782.000 ;
      RECT 635.400 18.000 639.000 782.000 ;
      RECT 664.200 18.000 667.800 782.000 ;
      RECT 693.000 18.000 696.600 782.000 ;
      RECT 721.800 18.000 725.400 782.000 ;
      RECT 750.600 18.000 754.200 782.000 ;
      RECT 779.400 18.000 783.000 782.000 ;
      RECT 808.200 18.000 811.800 782.000 ;
      RECT 837.000 18.000 840.600 782.000 ;
      RECT 865.800 18.000 869.400 782.000 ;
      RECT 894.600 18.000 898.200 782.000 ;
      RECT 923.400 18.000 927.000 782.000 ;
      RECT 952.200 18.000 955.800 782.000 ;
      RECT 981.000 18.000 984.600 782.000 ;
      RECT 1009.800 18.000 1013.400 782.000 ;
      RECT 1038.600 18.000 1042.200 782.000 ;
      RECT 1067.400 18.000 1071.000 782.000 ;
      RECT 1096.200 18.000 1099.800 782.000 ;
      RECT 1125.000 18.000 1128.600 782.000 ;
      RECT 1153.800 18.000 1157.400 782.000 ;
      RECT 1182.600 18.000 1186.200 782.000 ;
      RECT 1211.400 18.000 1215.000 782.000 ;
      RECT 1240.200 18.000 1243.800 782.000 ;
      RECT 1269.000 18.000 1272.600 782.000 ;
      RECT 1297.800 18.000 1301.400 782.000 ;
      RECT 1326.600 18.000 1330.200 782.000 ;
      RECT 1355.400 18.000 1359.000 782.000 ;
      RECT 1384.200 18.000 1387.800 782.000 ;
      RECT 1413.000 18.000 1416.600 782.000 ;
      RECT 1441.800 18.000 1445.400 782.000 ;
      RECT 1470.600 18.000 1474.200 782.000 ;
      RECT 1499.400 18.000 1503.000 782.000 ;
      RECT 1528.200 18.000 1531.800 782.000 ;
      RECT 1557.000 18.000 1560.600 782.000 ;
      RECT 1585.800 18.000 1589.400 782.000 ;
      RECT 1614.600 18.000 1618.200 782.000 ;
      RECT 1643.400 18.000 1647.000 782.000 ;
      RECT 1672.200 18.000 1675.800 782.000 ;
      RECT 1701.000 18.000 1704.600 782.000 ;
      RECT 1729.800 18.000 1733.400 782.000 ;
      RECT 1758.600 18.000 1762.200 782.000 ;
    END
  END vccd1
  OBS
    LAYER met1 ;
    RECT 0 0 1800.000 800.000 ;
    LAYER met2 ;
    RECT 0 0 1800.000 800.000 ;
    LAYER met3 ;
    RECT 0.900 0 1800.000 800.000 ;
    RECT 0 0.000 0.900 17.550 ;
    RECT 0 18.450 0.900 19.350 ;
    RECT 0 20.250 0.900 21.150 ;
    RECT 0 22.050 0.900 22.950 ;
    RECT 0 23.850 0.900 24.750 ;
    RECT 0 25.650 0.900 26.550 ;
    RECT 0 27.450 0.900 28.350 ;
    RECT 0 29.250 0.900 30.150 ;
    RECT 0 31.050 0.900 31.950 ;
    RECT 0 32.850 0.900 33.750 ;
    RECT 0 34.650 0.900 35.550 ;
    RECT 0 36.450 0.900 37.350 ;
    RECT 0 38.250 0.900 39.150 ;
    RECT 0 40.050 0.900 40.950 ;
    RECT 0 41.850 0.900 42.750 ;
    RECT 0 43.650 0.900 44.550 ;
    RECT 0 45.450 0.900 46.350 ;
    RECT 0 47.250 0.900 48.150 ;
    RECT 0 49.050 0.900 49.950 ;
    RECT 0 50.850 0.900 51.750 ;
    RECT 0 52.650 0.900 53.550 ;
    RECT 0 54.450 0.900 55.350 ;
    RECT 0 56.250 0.900 57.150 ;
    RECT 0 58.050 0.900 58.950 ;
    RECT 0 59.850 0.900 60.750 ;
    RECT 0 61.650 0.900 62.550 ;
    RECT 0 63.450 0.900 64.350 ;
    RECT 0 65.250 0.900 66.150 ;
    RECT 0 67.050 0.900 67.950 ;
    RECT 0 68.850 0.900 69.750 ;
    RECT 0 70.650 0.900 71.550 ;
    RECT 0 72.450 0.900 73.350 ;
    RECT 0 74.250 0.900 75.150 ;
    RECT 0 76.050 0.900 76.950 ;
    RECT 0 77.850 0.900 78.750 ;
    RECT 0 79.650 0.900 80.550 ;
    RECT 0 81.450 0.900 82.350 ;
    RECT 0 83.250 0.900 84.150 ;
    RECT 0 85.050 0.900 85.950 ;
    RECT 0 86.850 0.900 87.750 ;
    RECT 0 88.650 0.900 89.550 ;
    RECT 0 90.450 0.900 91.350 ;
    RECT 0 92.250 0.900 93.150 ;
    RECT 0 94.050 0.900 94.950 ;
    RECT 0 95.850 0.900 96.750 ;
    RECT 0 97.650 0.900 98.550 ;
    RECT 0 99.450 0.900 100.350 ;
    RECT 0 101.250 0.900 102.150 ;
    RECT 0 103.050 0.900 103.950 ;
    RECT 0 104.850 0.900 105.750 ;
    RECT 0 106.650 0.900 107.550 ;
    RECT 0 108.450 0.900 109.350 ;
    RECT 0 110.250 0.900 111.150 ;
    RECT 0 112.050 0.900 112.950 ;
    RECT 0 113.850 0.900 114.750 ;
    RECT 0 115.650 0.900 116.550 ;
    RECT 0 117.450 0.900 118.350 ;
    RECT 0 119.250 0.900 120.150 ;
    RECT 0 121.050 0.900 121.950 ;
    RECT 0 122.850 0.900 123.750 ;
    RECT 0 124.650 0.900 125.550 ;
    RECT 0 126.450 0.900 127.350 ;
    RECT 0 128.250 0.900 129.150 ;
    RECT 0 130.050 0.900 130.950 ;
    RECT 0 131.850 0.900 132.750 ;
    RECT 0 133.650 0.900 134.550 ;
    RECT 0 135.450 0.900 136.350 ;
    RECT 0 137.250 0.900 138.150 ;
    RECT 0 139.050 0.900 139.950 ;
    RECT 0 140.850 0.900 141.750 ;
    RECT 0 142.650 0.900 143.550 ;
    RECT 0 144.450 0.900 145.350 ;
    RECT 0 146.250 0.900 147.150 ;
    RECT 0 148.050 0.900 148.950 ;
    RECT 0 149.850 0.900 150.750 ;
    RECT 0 151.650 0.900 152.550 ;
    RECT 0 153.450 0.900 154.350 ;
    RECT 0 155.250 0.900 156.150 ;
    RECT 0 157.050 0.900 157.950 ;
    RECT 0 158.850 0.900 159.750 ;
    RECT 0 160.650 0.900 161.550 ;
    RECT 0 162.450 0.900 163.350 ;
    RECT 0 164.250 0.900 165.150 ;
    RECT 0 166.050 0.900 166.950 ;
    RECT 0 167.850 0.900 168.750 ;
    RECT 0 169.650 0.900 170.550 ;
    RECT 0 171.450 0.900 172.350 ;
    RECT 0 173.250 0.900 174.150 ;
    RECT 0 175.050 0.900 175.950 ;
    RECT 0 176.850 0.900 177.750 ;
    RECT 0 178.650 0.900 179.550 ;
    RECT 0 180.450 0.900 181.350 ;
    RECT 0 182.250 0.900 183.150 ;
    RECT 0 184.050 0.900 184.950 ;
    RECT 0 185.850 0.900 186.750 ;
    RECT 0 187.650 0.900 188.550 ;
    RECT 0 189.450 0.900 244.350 ;
    RECT 0 245.250 0.900 246.150 ;
    RECT 0 247.050 0.900 247.950 ;
    RECT 0 248.850 0.900 249.750 ;
    RECT 0 250.650 0.900 251.550 ;
    RECT 0 252.450 0.900 253.350 ;
    RECT 0 254.250 0.900 255.150 ;
    RECT 0 256.050 0.900 256.950 ;
    RECT 0 257.850 0.900 258.750 ;
    RECT 0 259.650 0.900 260.550 ;
    RECT 0 261.450 0.900 262.350 ;
    RECT 0 263.250 0.900 264.150 ;
    RECT 0 265.050 0.900 265.950 ;
    RECT 0 266.850 0.900 267.750 ;
    RECT 0 268.650 0.900 269.550 ;
    RECT 0 270.450 0.900 271.350 ;
    RECT 0 272.250 0.900 273.150 ;
    RECT 0 274.050 0.900 274.950 ;
    RECT 0 275.850 0.900 276.750 ;
    RECT 0 277.650 0.900 278.550 ;
    RECT 0 279.450 0.900 280.350 ;
    RECT 0 281.250 0.900 282.150 ;
    RECT 0 283.050 0.900 283.950 ;
    RECT 0 284.850 0.900 285.750 ;
    RECT 0 286.650 0.900 287.550 ;
    RECT 0 288.450 0.900 289.350 ;
    RECT 0 290.250 0.900 291.150 ;
    RECT 0 292.050 0.900 292.950 ;
    RECT 0 293.850 0.900 294.750 ;
    RECT 0 295.650 0.900 296.550 ;
    RECT 0 297.450 0.900 298.350 ;
    RECT 0 299.250 0.900 300.150 ;
    RECT 0 301.050 0.900 301.950 ;
    RECT 0 302.850 0.900 303.750 ;
    RECT 0 304.650 0.900 305.550 ;
    RECT 0 306.450 0.900 307.350 ;
    RECT 0 308.250 0.900 309.150 ;
    RECT 0 310.050 0.900 310.950 ;
    RECT 0 311.850 0.900 312.750 ;
    RECT 0 313.650 0.900 314.550 ;
    RECT 0 315.450 0.900 316.350 ;
    RECT 0 317.250 0.900 318.150 ;
    RECT 0 319.050 0.900 319.950 ;
    RECT 0 320.850 0.900 321.750 ;
    RECT 0 322.650 0.900 323.550 ;
    RECT 0 324.450 0.900 325.350 ;
    RECT 0 326.250 0.900 327.150 ;
    RECT 0 328.050 0.900 328.950 ;
    RECT 0 329.850 0.900 330.750 ;
    RECT 0 331.650 0.900 332.550 ;
    RECT 0 333.450 0.900 334.350 ;
    RECT 0 335.250 0.900 336.150 ;
    RECT 0 337.050 0.900 337.950 ;
    RECT 0 338.850 0.900 339.750 ;
    RECT 0 340.650 0.900 341.550 ;
    RECT 0 342.450 0.900 343.350 ;
    RECT 0 344.250 0.900 345.150 ;
    RECT 0 346.050 0.900 346.950 ;
    RECT 0 347.850 0.900 348.750 ;
    RECT 0 349.650 0.900 350.550 ;
    RECT 0 351.450 0.900 352.350 ;
    RECT 0 353.250 0.900 354.150 ;
    RECT 0 355.050 0.900 355.950 ;
    RECT 0 356.850 0.900 357.750 ;
    RECT 0 358.650 0.900 359.550 ;
    RECT 0 360.450 0.900 361.350 ;
    RECT 0 362.250 0.900 363.150 ;
    RECT 0 364.050 0.900 364.950 ;
    RECT 0 365.850 0.900 366.750 ;
    RECT 0 367.650 0.900 368.550 ;
    RECT 0 369.450 0.900 370.350 ;
    RECT 0 371.250 0.900 372.150 ;
    RECT 0 373.050 0.900 373.950 ;
    RECT 0 374.850 0.900 375.750 ;
    RECT 0 376.650 0.900 377.550 ;
    RECT 0 378.450 0.900 379.350 ;
    RECT 0 380.250 0.900 381.150 ;
    RECT 0 382.050 0.900 382.950 ;
    RECT 0 383.850 0.900 384.750 ;
    RECT 0 385.650 0.900 386.550 ;
    RECT 0 387.450 0.900 388.350 ;
    RECT 0 389.250 0.900 390.150 ;
    RECT 0 391.050 0.900 391.950 ;
    RECT 0 392.850 0.900 393.750 ;
    RECT 0 394.650 0.900 395.550 ;
    RECT 0 396.450 0.900 397.350 ;
    RECT 0 398.250 0.900 399.150 ;
    RECT 0 400.050 0.900 400.950 ;
    RECT 0 401.850 0.900 402.750 ;
    RECT 0 403.650 0.900 404.550 ;
    RECT 0 405.450 0.900 406.350 ;
    RECT 0 407.250 0.900 408.150 ;
    RECT 0 409.050 0.900 409.950 ;
    RECT 0 410.850 0.900 411.750 ;
    RECT 0 412.650 0.900 413.550 ;
    RECT 0 414.450 0.900 415.350 ;
    RECT 0 416.250 0.900 471.150 ;
    RECT 0 472.050 0.900 472.950 ;
    RECT 0 473.850 0.900 474.750 ;
    RECT 0 475.650 0.900 476.550 ;
    RECT 0 477.450 0.900 478.350 ;
    RECT 0 479.250 0.900 480.150 ;
    RECT 0 481.050 0.900 481.950 ;
    RECT 0 482.850 0.900 483.750 ;
    RECT 0 484.650 0.900 485.550 ;
    RECT 0 486.450 0.900 487.350 ;
    RECT 0 488.250 0.900 489.150 ;
    RECT 0 490.050 0.900 490.950 ;
    RECT 0 491.850 0.900 492.750 ;
    RECT 0 493.650 0.900 494.550 ;
    RECT 0 495.450 0.900 496.350 ;
    RECT 0 497.250 0.900 498.150 ;
    RECT 0 499.050 0.900 499.950 ;
    RECT 0 500.850 0.900 501.750 ;
    RECT 0 502.650 0.900 503.550 ;
    RECT 0 504.450 0.900 505.350 ;
    RECT 0 506.250 0.900 507.150 ;
    RECT 0 508.050 0.900 508.950 ;
    RECT 0 509.850 0.900 510.750 ;
    RECT 0 511.650 0.900 512.550 ;
    RECT 0 513.450 0.900 514.350 ;
    RECT 0 515.250 0.900 516.150 ;
    RECT 0 517.050 0.900 517.950 ;
    RECT 0 518.850 0.900 519.750 ;
    RECT 0 520.650 0.900 521.550 ;
    RECT 0 522.450 0.900 523.350 ;
    RECT 0 524.250 0.900 525.150 ;
    RECT 0 526.050 0.900 526.950 ;
    RECT 0 527.850 0.900 528.750 ;
    RECT 0 529.650 0.900 530.550 ;
    RECT 0 531.450 0.900 532.350 ;
    RECT 0 533.250 0.900 534.150 ;
    RECT 0 535.050 0.900 535.950 ;
    RECT 0 536.850 0.900 537.750 ;
    RECT 0 538.650 0.900 539.550 ;
    RECT 0 540.450 0.900 541.350 ;
    RECT 0 542.250 0.900 543.150 ;
    RECT 0 544.050 0.900 544.950 ;
    RECT 0 545.850 0.900 546.750 ;
    RECT 0 547.650 0.900 548.550 ;
    RECT 0 549.450 0.900 550.350 ;
    RECT 0 551.250 0.900 552.150 ;
    RECT 0 553.050 0.900 553.950 ;
    RECT 0 554.850 0.900 555.750 ;
    RECT 0 556.650 0.900 557.550 ;
    RECT 0 558.450 0.900 559.350 ;
    RECT 0 560.250 0.900 561.150 ;
    RECT 0 562.050 0.900 562.950 ;
    RECT 0 563.850 0.900 564.750 ;
    RECT 0 565.650 0.900 566.550 ;
    RECT 0 567.450 0.900 568.350 ;
    RECT 0 569.250 0.900 570.150 ;
    RECT 0 571.050 0.900 571.950 ;
    RECT 0 572.850 0.900 573.750 ;
    RECT 0 574.650 0.900 575.550 ;
    RECT 0 576.450 0.900 577.350 ;
    RECT 0 578.250 0.900 579.150 ;
    RECT 0 580.050 0.900 580.950 ;
    RECT 0 581.850 0.900 582.750 ;
    RECT 0 583.650 0.900 584.550 ;
    RECT 0 585.450 0.900 586.350 ;
    RECT 0 587.250 0.900 588.150 ;
    RECT 0 589.050 0.900 589.950 ;
    RECT 0 590.850 0.900 591.750 ;
    RECT 0 592.650 0.900 593.550 ;
    RECT 0 594.450 0.900 595.350 ;
    RECT 0 596.250 0.900 597.150 ;
    RECT 0 598.050 0.900 598.950 ;
    RECT 0 599.850 0.900 600.750 ;
    RECT 0 601.650 0.900 602.550 ;
    RECT 0 603.450 0.900 604.350 ;
    RECT 0 605.250 0.900 606.150 ;
    RECT 0 607.050 0.900 607.950 ;
    RECT 0 608.850 0.900 609.750 ;
    RECT 0 610.650 0.900 611.550 ;
    RECT 0 612.450 0.900 613.350 ;
    RECT 0 614.250 0.900 615.150 ;
    RECT 0 616.050 0.900 616.950 ;
    RECT 0 617.850 0.900 618.750 ;
    RECT 0 619.650 0.900 620.550 ;
    RECT 0 621.450 0.900 622.350 ;
    RECT 0 623.250 0.900 624.150 ;
    RECT 0 625.050 0.900 625.950 ;
    RECT 0 626.850 0.900 627.750 ;
    RECT 0 628.650 0.900 629.550 ;
    RECT 0 630.450 0.900 631.350 ;
    RECT 0 632.250 0.900 633.150 ;
    RECT 0 634.050 0.900 634.950 ;
    RECT 0 635.850 0.900 636.750 ;
    RECT 0 637.650 0.900 638.550 ;
    RECT 0 639.450 0.900 640.350 ;
    RECT 0 641.250 0.900 642.150 ;
    RECT 0 643.050 0.900 697.950 ;
    RECT 0 698.850 0.900 699.750 ;
    RECT 0 700.650 0.900 701.550 ;
    RECT 0 702.450 0.900 703.350 ;
    RECT 0 704.250 0.900 705.150 ;
    RECT 0 706.050 0.900 706.950 ;
    RECT 0 707.850 0.900 762.750 ;
    RECT 0 763.650 0.900 764.550 ;
    RECT 0 765.450 0.900 766.350 ;
    RECT 0 767.250 0.900 800.000 ;
    LAYER met4 ;
    RECT 0 0 1800.000 18.000 ;
    RECT 0 782.000 1800.000 800.000 ;
    RECT 0.000 18.000 16.200 782.000 ;
    RECT 19.800 18.000 30.600 782.000 ;
    RECT 34.200 18.000 45.000 782.000 ;
    RECT 48.600 18.000 59.400 782.000 ;
    RECT 63.000 18.000 73.800 782.000 ;
    RECT 77.400 18.000 88.200 782.000 ;
    RECT 91.800 18.000 102.600 782.000 ;
    RECT 106.200 18.000 117.000 782.000 ;
    RECT 120.600 18.000 131.400 782.000 ;
    RECT 135.000 18.000 145.800 782.000 ;
    RECT 149.400 18.000 160.200 782.000 ;
    RECT 163.800 18.000 174.600 782.000 ;
    RECT 178.200 18.000 189.000 782.000 ;
    RECT 192.600 18.000 203.400 782.000 ;
    RECT 207.000 18.000 217.800 782.000 ;
    RECT 221.400 18.000 232.200 782.000 ;
    RECT 235.800 18.000 246.600 782.000 ;
    RECT 250.200 18.000 261.000 782.000 ;
    RECT 264.600 18.000 275.400 782.000 ;
    RECT 279.000 18.000 289.800 782.000 ;
    RECT 293.400 18.000 304.200 782.000 ;
    RECT 307.800 18.000 318.600 782.000 ;
    RECT 322.200 18.000 333.000 782.000 ;
    RECT 336.600 18.000 347.400 782.000 ;
    RECT 351.000 18.000 361.800 782.000 ;
    RECT 365.400 18.000 376.200 782.000 ;
    RECT 379.800 18.000 390.600 782.000 ;
    RECT 394.200 18.000 405.000 782.000 ;
    RECT 408.600 18.000 419.400 782.000 ;
    RECT 423.000 18.000 433.800 782.000 ;
    RECT 437.400 18.000 448.200 782.000 ;
    RECT 451.800 18.000 462.600 782.000 ;
    RECT 466.200 18.000 477.000 782.000 ;
    RECT 480.600 18.000 491.400 782.000 ;
    RECT 495.000 18.000 505.800 782.000 ;
    RECT 509.400 18.000 520.200 782.000 ;
    RECT 523.800 18.000 534.600 782.000 ;
    RECT 538.200 18.000 549.000 782.000 ;
    RECT 552.600 18.000 563.400 782.000 ;
    RECT 567.000 18.000 577.800 782.000 ;
    RECT 581.400 18.000 592.200 782.000 ;
    RECT 595.800 18.000 606.600 782.000 ;
    RECT 610.200 18.000 621.000 782.000 ;
    RECT 624.600 18.000 635.400 782.000 ;
    RECT 639.000 18.000 649.800 782.000 ;
    RECT 653.400 18.000 664.200 782.000 ;
    RECT 667.800 18.000 678.600 782.000 ;
    RECT 682.200 18.000 693.000 782.000 ;
    RECT 696.600 18.000 707.400 782.000 ;
    RECT 711.000 18.000 721.800 782.000 ;
    RECT 725.400 18.000 736.200 782.000 ;
    RECT 739.800 18.000 750.600 782.000 ;
    RECT 754.200 18.000 765.000 782.000 ;
    RECT 768.600 18.000 779.400 782.000 ;
    RECT 783.000 18.000 793.800 782.000 ;
    RECT 797.400 18.000 808.200 782.000 ;
    RECT 811.800 18.000 822.600 782.000 ;
    RECT 826.200 18.000 837.000 782.000 ;
    RECT 840.600 18.000 851.400 782.000 ;
    RECT 855.000 18.000 865.800 782.000 ;
    RECT 869.400 18.000 880.200 782.000 ;
    RECT 883.800 18.000 894.600 782.000 ;
    RECT 898.200 18.000 909.000 782.000 ;
    RECT 912.600 18.000 923.400 782.000 ;
    RECT 927.000 18.000 937.800 782.000 ;
    RECT 941.400 18.000 952.200 782.000 ;
    RECT 955.800 18.000 966.600 782.000 ;
    RECT 970.200 18.000 981.000 782.000 ;
    RECT 984.600 18.000 995.400 782.000 ;
    RECT 999.000 18.000 1009.800 782.000 ;
    RECT 1013.400 18.000 1024.200 782.000 ;
    RECT 1027.800 18.000 1038.600 782.000 ;
    RECT 1042.200 18.000 1053.000 782.000 ;
    RECT 1056.600 18.000 1067.400 782.000 ;
    RECT 1071.000 18.000 1081.800 782.000 ;
    RECT 1085.400 18.000 1096.200 782.000 ;
    RECT 1099.800 18.000 1110.600 782.000 ;
    RECT 1114.200 18.000 1125.000 782.000 ;
    RECT 1128.600 18.000 1139.400 782.000 ;
    RECT 1143.000 18.000 1153.800 782.000 ;
    RECT 1157.400 18.000 1168.200 782.000 ;
    RECT 1171.800 18.000 1182.600 782.000 ;
    RECT 1186.200 18.000 1197.000 782.000 ;
    RECT 1200.600 18.000 1211.400 782.000 ;
    RECT 1215.000 18.000 1225.800 782.000 ;
    RECT 1229.400 18.000 1240.200 782.000 ;
    RECT 1243.800 18.000 1254.600 782.000 ;
    RECT 1258.200 18.000 1269.000 782.000 ;
    RECT 1272.600 18.000 1283.400 782.000 ;
    RECT 1287.000 18.000 1297.800 782.000 ;
    RECT 1301.400 18.000 1312.200 782.000 ;
    RECT 1315.800 18.000 1326.600 782.000 ;
    RECT 1330.200 18.000 1341.000 782.000 ;
    RECT 1344.600 18.000 1355.400 782.000 ;
    RECT 1359.000 18.000 1369.800 782.000 ;
    RECT 1373.400 18.000 1384.200 782.000 ;
    RECT 1387.800 18.000 1398.600 782.000 ;
    RECT 1402.200 18.000 1413.000 782.000 ;
    RECT 1416.600 18.000 1427.400 782.000 ;
    RECT 1431.000 18.000 1441.800 782.000 ;
    RECT 1445.400 18.000 1456.200 782.000 ;
    RECT 1459.800 18.000 1470.600 782.000 ;
    RECT 1474.200 18.000 1485.000 782.000 ;
    RECT 1488.600 18.000 1499.400 782.000 ;
    RECT 1503.000 18.000 1513.800 782.000 ;
    RECT 1517.400 18.000 1528.200 782.000 ;
    RECT 1531.800 18.000 1542.600 782.000 ;
    RECT 1546.200 18.000 1557.000 782.000 ;
    RECT 1560.600 18.000 1571.400 782.000 ;
    RECT 1575.000 18.000 1585.800 782.000 ;
    RECT 1589.400 18.000 1600.200 782.000 ;
    RECT 1603.800 18.000 1614.600 782.000 ;
    RECT 1618.200 18.000 1629.000 782.000 ;
    RECT 1632.600 18.000 1643.400 782.000 ;
    RECT 1647.000 18.000 1657.800 782.000 ;
    RECT 1661.400 18.000 1672.200 782.000 ;
    RECT 1675.800 18.000 1686.600 782.000 ;
    RECT 1690.200 18.000 1701.000 782.000 ;
    RECT 1704.600 18.000 1715.400 782.000 ;
    RECT 1719.000 18.000 1729.800 782.000 ;
    RECT 1733.400 18.000 1744.200 782.000 ;
    RECT 1747.800 18.000 1758.600 782.000 ;
    RECT 1762.200 18.000 1773.000 782.000 ;
    RECT 1776.600 18.000 1800.000 782.000 ;

  END
END fakeram130_64x96

END LIBRARY
