VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_512x64
  FOREIGN fakeram130_512x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 316.800 BY 657.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.200 0.600 6.800 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.800 0.600 9.400 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 11.400 0.600 12.000 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.000 0.600 14.600 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.600 0.600 17.200 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 19.200 0.600 19.800 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.800 0.600 22.400 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.400 0.600 25.000 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.000 0.600 27.600 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.600 0.600 30.200 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.200 0.600 32.800 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.800 0.600 35.400 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.400 0.600 38.000 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.000 0.600 40.600 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.600 0.600 43.200 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.200 0.600 45.800 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.800 0.600 48.400 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.400 0.600 51.000 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 53.000 0.600 53.600 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.600 0.600 56.200 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 58.200 0.600 58.800 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 60.800 0.600 61.400 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.400 0.600 64.000 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.000 0.600 66.600 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 68.600 0.600 69.200 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.200 0.600 71.800 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.800 0.600 74.400 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.400 0.600 77.000 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.000 0.600 79.600 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.600 0.600 82.200 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.200 0.600 84.800 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.800 0.600 87.400 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.400 0.600 90.000 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.000 0.600 92.600 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.600 0.600 95.200 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.200 0.600 97.800 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.800 0.600 100.400 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.400 0.600 103.000 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.000 0.600 105.600 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 107.600 0.600 108.200 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.200 0.600 110.800 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 112.800 0.600 113.400 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 115.400 0.600 116.000 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.000 0.600 118.600 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 120.600 0.600 121.200 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 123.200 0.600 123.800 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 125.800 0.600 126.400 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 128.400 0.600 129.000 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.000 0.600 131.600 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.600 0.600 134.200 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.200 0.600 136.800 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 138.800 0.600 139.400 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.400 0.600 142.000 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.000 0.600 144.600 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.600 0.600 147.200 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.200 0.600 149.800 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.800 0.600 152.400 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.400 0.600 155.000 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.000 0.600 157.600 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 159.600 0.600 160.200 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.200 0.600 162.800 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.800 0.600 165.400 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.400 0.600 168.000 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 170.000 0.600 170.600 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 197.950 0.600 198.550 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 200.550 0.600 201.150 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 203.150 0.600 203.750 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.750 0.600 206.350 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 208.350 0.600 208.950 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 210.950 0.600 211.550 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 213.550 0.600 214.150 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.150 0.600 216.750 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 218.750 0.600 219.350 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 221.350 0.600 221.950 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.950 0.600 224.550 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 226.550 0.600 227.150 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 229.150 0.600 229.750 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 231.750 0.600 232.350 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 234.350 0.600 234.950 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 236.950 0.600 237.550 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 239.550 0.600 240.150 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 242.150 0.600 242.750 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 244.750 0.600 245.350 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 247.350 0.600 247.950 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 249.950 0.600 250.550 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 252.550 0.600 253.150 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 255.150 0.600 255.750 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 257.750 0.600 258.350 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 260.350 0.600 260.950 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 262.950 0.600 263.550 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 265.550 0.600 266.150 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 268.150 0.600 268.750 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 270.750 0.600 271.350 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 273.350 0.600 273.950 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 275.950 0.600 276.550 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 278.550 0.600 279.150 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 281.150 0.600 281.750 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 283.750 0.600 284.350 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 286.350 0.600 286.950 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 288.950 0.600 289.550 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 291.550 0.600 292.150 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 294.150 0.600 294.750 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 296.750 0.600 297.350 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 299.350 0.600 299.950 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 301.950 0.600 302.550 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 304.550 0.600 305.150 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 307.150 0.600 307.750 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 309.750 0.600 310.350 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 312.350 0.600 312.950 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 314.950 0.600 315.550 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 317.550 0.600 318.150 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 320.150 0.600 320.750 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 322.750 0.600 323.350 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 325.350 0.600 325.950 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.950 0.600 328.550 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 330.550 0.600 331.150 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.150 0.600 333.750 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 335.750 0.600 336.350 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 338.350 0.600 338.950 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 340.950 0.600 341.550 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 343.550 0.600 344.150 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 346.150 0.600 346.750 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 348.750 0.600 349.350 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 351.350 0.600 351.950 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 353.950 0.600 354.550 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 356.550 0.600 357.150 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 359.150 0.600 359.750 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 361.750 0.600 362.350 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 389.700 0.600 390.300 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 392.300 0.600 392.900 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 394.900 0.600 395.500 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 397.500 0.600 398.100 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 400.100 0.600 400.700 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 402.700 0.600 403.300 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 405.300 0.600 405.900 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 407.900 0.600 408.500 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 410.500 0.600 411.100 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 413.100 0.600 413.700 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 415.700 0.600 416.300 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 418.300 0.600 418.900 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 420.900 0.600 421.500 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 423.500 0.600 424.100 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 426.100 0.600 426.700 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 428.700 0.600 429.300 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 431.300 0.600 431.900 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 433.900 0.600 434.500 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 436.500 0.600 437.100 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 439.100 0.600 439.700 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 441.700 0.600 442.300 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 444.300 0.600 444.900 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 446.900 0.600 447.500 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 449.500 0.600 450.100 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 452.100 0.600 452.700 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 454.700 0.600 455.300 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 457.300 0.600 457.900 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 459.900 0.600 460.500 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 462.500 0.600 463.100 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 465.100 0.600 465.700 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 467.700 0.600 468.300 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 470.300 0.600 470.900 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 472.900 0.600 473.500 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 475.500 0.600 476.100 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 478.100 0.600 478.700 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 480.700 0.600 481.300 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 483.300 0.600 483.900 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.900 0.600 486.500 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 488.500 0.600 489.100 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 491.100 0.600 491.700 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 493.700 0.600 494.300 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 496.300 0.600 496.900 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 498.900 0.600 499.500 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.500 0.600 502.100 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 504.100 0.600 504.700 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 506.700 0.600 507.300 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 509.300 0.600 509.900 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 511.900 0.600 512.500 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 514.500 0.600 515.100 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 517.100 0.600 517.700 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 519.700 0.600 520.300 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 522.300 0.600 522.900 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 524.900 0.600 525.500 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 527.500 0.600 528.100 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 530.100 0.600 530.700 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 532.700 0.600 533.300 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.300 0.600 535.900 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 537.900 0.600 538.500 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 540.500 0.600 541.100 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 543.100 0.600 543.700 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 545.700 0.600 546.300 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 548.300 0.600 548.900 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 550.900 0.600 551.500 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 553.500 0.600 554.100 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 581.450 0.600 582.050 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 584.050 0.600 584.650 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 586.650 0.600 587.250 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 589.250 0.600 589.850 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 591.850 0.600 592.450 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 594.450 0.600 595.050 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 597.050 0.600 597.650 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 599.650 0.600 600.250 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 602.250 0.600 602.850 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 630.200 0.600 630.800 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 632.800 0.600 633.400 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 635.400 0.600 636.000 ;
    END
  END clk
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 5.300 6.500 7.700 650.500 ;
      RECT 15.700 6.500 18.100 650.500 ;
      RECT 26.100 6.500 28.500 650.500 ;
      RECT 36.500 6.500 38.900 650.500 ;
      RECT 46.900 6.500 49.300 650.500 ;
      RECT 57.300 6.500 59.700 650.500 ;
      RECT 67.700 6.500 70.100 650.500 ;
      RECT 78.100 6.500 80.500 650.500 ;
      RECT 88.500 6.500 90.900 650.500 ;
      RECT 98.900 6.500 101.300 650.500 ;
      RECT 109.300 6.500 111.700 650.500 ;
      RECT 119.700 6.500 122.100 650.500 ;
      RECT 130.100 6.500 132.500 650.500 ;
      RECT 140.500 6.500 142.900 650.500 ;
      RECT 150.900 6.500 153.300 650.500 ;
      RECT 161.300 6.500 163.700 650.500 ;
      RECT 171.700 6.500 174.100 650.500 ;
      RECT 182.100 6.500 184.500 650.500 ;
      RECT 192.500 6.500 194.900 650.500 ;
      RECT 202.900 6.500 205.300 650.500 ;
      RECT 213.300 6.500 215.700 650.500 ;
      RECT 223.700 6.500 226.100 650.500 ;
      RECT 234.100 6.500 236.500 650.500 ;
      RECT 244.500 6.500 246.900 650.500 ;
      RECT 254.900 6.500 257.300 650.500 ;
      RECT 265.300 6.500 267.700 650.500 ;
      RECT 275.700 6.500 278.100 650.500 ;
      RECT 286.100 6.500 288.500 650.500 ;
      RECT 296.500 6.500 298.900 650.500 ;
      RECT 306.900 6.500 309.300 650.500 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 10.500 6.500 12.900 650.500 ;
      RECT 20.900 6.500 23.300 650.500 ;
      RECT 31.300 6.500 33.700 650.500 ;
      RECT 41.700 6.500 44.100 650.500 ;
      RECT 52.100 6.500 54.500 650.500 ;
      RECT 62.500 6.500 64.900 650.500 ;
      RECT 72.900 6.500 75.300 650.500 ;
      RECT 83.300 6.500 85.700 650.500 ;
      RECT 93.700 6.500 96.100 650.500 ;
      RECT 104.100 6.500 106.500 650.500 ;
      RECT 114.500 6.500 116.900 650.500 ;
      RECT 124.900 6.500 127.300 650.500 ;
      RECT 135.300 6.500 137.700 650.500 ;
      RECT 145.700 6.500 148.100 650.500 ;
      RECT 156.100 6.500 158.500 650.500 ;
      RECT 166.500 6.500 168.900 650.500 ;
      RECT 176.900 6.500 179.300 650.500 ;
      RECT 187.300 6.500 189.700 650.500 ;
      RECT 197.700 6.500 200.100 650.500 ;
      RECT 208.100 6.500 210.500 650.500 ;
      RECT 218.500 6.500 220.900 650.500 ;
      RECT 228.900 6.500 231.300 650.500 ;
      RECT 239.300 6.500 241.700 650.500 ;
      RECT 249.700 6.500 252.100 650.500 ;
      RECT 260.100 6.500 262.500 650.500 ;
      RECT 270.500 6.500 272.900 650.500 ;
      RECT 280.900 6.500 283.300 650.500 ;
      RECT 291.300 6.500 293.700 650.500 ;
      RECT 301.700 6.500 304.100 650.500 ;
    END
  END VPWR
  OBS
    LAYER met1 ;
    RECT 0 0 316.800 657.000 ;
    LAYER met2 ;
    RECT 0 0 316.800 657.000 ;
    LAYER met3 ;
    RECT 0.600 0 316.800 657.000 ;
    RECT 0 0.000 0.600 6.200 ;
    RECT 0 6.800 0.600 8.800 ;
    RECT 0 9.400 0.600 11.400 ;
    RECT 0 12.000 0.600 14.000 ;
    RECT 0 14.600 0.600 16.600 ;
    RECT 0 17.200 0.600 19.200 ;
    RECT 0 19.800 0.600 21.800 ;
    RECT 0 22.400 0.600 24.400 ;
    RECT 0 25.000 0.600 27.000 ;
    RECT 0 27.600 0.600 29.600 ;
    RECT 0 30.200 0.600 32.200 ;
    RECT 0 32.800 0.600 34.800 ;
    RECT 0 35.400 0.600 37.400 ;
    RECT 0 38.000 0.600 40.000 ;
    RECT 0 40.600 0.600 42.600 ;
    RECT 0 43.200 0.600 45.200 ;
    RECT 0 45.800 0.600 47.800 ;
    RECT 0 48.400 0.600 50.400 ;
    RECT 0 51.000 0.600 53.000 ;
    RECT 0 53.600 0.600 55.600 ;
    RECT 0 56.200 0.600 58.200 ;
    RECT 0 58.800 0.600 60.800 ;
    RECT 0 61.400 0.600 63.400 ;
    RECT 0 64.000 0.600 66.000 ;
    RECT 0 66.600 0.600 68.600 ;
    RECT 0 69.200 0.600 71.200 ;
    RECT 0 71.800 0.600 73.800 ;
    RECT 0 74.400 0.600 76.400 ;
    RECT 0 77.000 0.600 79.000 ;
    RECT 0 79.600 0.600 81.600 ;
    RECT 0 82.200 0.600 84.200 ;
    RECT 0 84.800 0.600 86.800 ;
    RECT 0 87.400 0.600 89.400 ;
    RECT 0 90.000 0.600 92.000 ;
    RECT 0 92.600 0.600 94.600 ;
    RECT 0 95.200 0.600 97.200 ;
    RECT 0 97.800 0.600 99.800 ;
    RECT 0 100.400 0.600 102.400 ;
    RECT 0 103.000 0.600 105.000 ;
    RECT 0 105.600 0.600 107.600 ;
    RECT 0 108.200 0.600 110.200 ;
    RECT 0 110.800 0.600 112.800 ;
    RECT 0 113.400 0.600 115.400 ;
    RECT 0 116.000 0.600 118.000 ;
    RECT 0 118.600 0.600 120.600 ;
    RECT 0 121.200 0.600 123.200 ;
    RECT 0 123.800 0.600 125.800 ;
    RECT 0 126.400 0.600 128.400 ;
    RECT 0 129.000 0.600 131.000 ;
    RECT 0 131.600 0.600 133.600 ;
    RECT 0 134.200 0.600 136.200 ;
    RECT 0 136.800 0.600 138.800 ;
    RECT 0 139.400 0.600 141.400 ;
    RECT 0 142.000 0.600 144.000 ;
    RECT 0 144.600 0.600 146.600 ;
    RECT 0 147.200 0.600 149.200 ;
    RECT 0 149.800 0.600 151.800 ;
    RECT 0 152.400 0.600 154.400 ;
    RECT 0 155.000 0.600 157.000 ;
    RECT 0 157.600 0.600 159.600 ;
    RECT 0 160.200 0.600 162.200 ;
    RECT 0 162.800 0.600 164.800 ;
    RECT 0 165.400 0.600 167.400 ;
    RECT 0 168.000 0.600 170.000 ;
    RECT 0 170.600 0.600 197.950 ;
    RECT 0 198.550 0.600 200.550 ;
    RECT 0 201.150 0.600 203.150 ;
    RECT 0 203.750 0.600 205.750 ;
    RECT 0 206.350 0.600 208.350 ;
    RECT 0 208.950 0.600 210.950 ;
    RECT 0 211.550 0.600 213.550 ;
    RECT 0 214.150 0.600 216.150 ;
    RECT 0 216.750 0.600 218.750 ;
    RECT 0 219.350 0.600 221.350 ;
    RECT 0 221.950 0.600 223.950 ;
    RECT 0 224.550 0.600 226.550 ;
    RECT 0 227.150 0.600 229.150 ;
    RECT 0 229.750 0.600 231.750 ;
    RECT 0 232.350 0.600 234.350 ;
    RECT 0 234.950 0.600 236.950 ;
    RECT 0 237.550 0.600 239.550 ;
    RECT 0 240.150 0.600 242.150 ;
    RECT 0 242.750 0.600 244.750 ;
    RECT 0 245.350 0.600 247.350 ;
    RECT 0 247.950 0.600 249.950 ;
    RECT 0 250.550 0.600 252.550 ;
    RECT 0 253.150 0.600 255.150 ;
    RECT 0 255.750 0.600 257.750 ;
    RECT 0 258.350 0.600 260.350 ;
    RECT 0 260.950 0.600 262.950 ;
    RECT 0 263.550 0.600 265.550 ;
    RECT 0 266.150 0.600 268.150 ;
    RECT 0 268.750 0.600 270.750 ;
    RECT 0 271.350 0.600 273.350 ;
    RECT 0 273.950 0.600 275.950 ;
    RECT 0 276.550 0.600 278.550 ;
    RECT 0 279.150 0.600 281.150 ;
    RECT 0 281.750 0.600 283.750 ;
    RECT 0 284.350 0.600 286.350 ;
    RECT 0 286.950 0.600 288.950 ;
    RECT 0 289.550 0.600 291.550 ;
    RECT 0 292.150 0.600 294.150 ;
    RECT 0 294.750 0.600 296.750 ;
    RECT 0 297.350 0.600 299.350 ;
    RECT 0 299.950 0.600 301.950 ;
    RECT 0 302.550 0.600 304.550 ;
    RECT 0 305.150 0.600 307.150 ;
    RECT 0 307.750 0.600 309.750 ;
    RECT 0 310.350 0.600 312.350 ;
    RECT 0 312.950 0.600 314.950 ;
    RECT 0 315.550 0.600 317.550 ;
    RECT 0 318.150 0.600 320.150 ;
    RECT 0 320.750 0.600 322.750 ;
    RECT 0 323.350 0.600 325.350 ;
    RECT 0 325.950 0.600 327.950 ;
    RECT 0 328.550 0.600 330.550 ;
    RECT 0 331.150 0.600 333.150 ;
    RECT 0 333.750 0.600 335.750 ;
    RECT 0 336.350 0.600 338.350 ;
    RECT 0 338.950 0.600 340.950 ;
    RECT 0 341.550 0.600 343.550 ;
    RECT 0 344.150 0.600 346.150 ;
    RECT 0 346.750 0.600 348.750 ;
    RECT 0 349.350 0.600 351.350 ;
    RECT 0 351.950 0.600 353.950 ;
    RECT 0 354.550 0.600 356.550 ;
    RECT 0 357.150 0.600 359.150 ;
    RECT 0 359.750 0.600 361.750 ;
    RECT 0 362.350 0.600 389.700 ;
    RECT 0 390.300 0.600 392.300 ;
    RECT 0 392.900 0.600 394.900 ;
    RECT 0 395.500 0.600 397.500 ;
    RECT 0 398.100 0.600 400.100 ;
    RECT 0 400.700 0.600 402.700 ;
    RECT 0 403.300 0.600 405.300 ;
    RECT 0 405.900 0.600 407.900 ;
    RECT 0 408.500 0.600 410.500 ;
    RECT 0 411.100 0.600 413.100 ;
    RECT 0 413.700 0.600 415.700 ;
    RECT 0 416.300 0.600 418.300 ;
    RECT 0 418.900 0.600 420.900 ;
    RECT 0 421.500 0.600 423.500 ;
    RECT 0 424.100 0.600 426.100 ;
    RECT 0 426.700 0.600 428.700 ;
    RECT 0 429.300 0.600 431.300 ;
    RECT 0 431.900 0.600 433.900 ;
    RECT 0 434.500 0.600 436.500 ;
    RECT 0 437.100 0.600 439.100 ;
    RECT 0 439.700 0.600 441.700 ;
    RECT 0 442.300 0.600 444.300 ;
    RECT 0 444.900 0.600 446.900 ;
    RECT 0 447.500 0.600 449.500 ;
    RECT 0 450.100 0.600 452.100 ;
    RECT 0 452.700 0.600 454.700 ;
    RECT 0 455.300 0.600 457.300 ;
    RECT 0 457.900 0.600 459.900 ;
    RECT 0 460.500 0.600 462.500 ;
    RECT 0 463.100 0.600 465.100 ;
    RECT 0 465.700 0.600 467.700 ;
    RECT 0 468.300 0.600 470.300 ;
    RECT 0 470.900 0.600 472.900 ;
    RECT 0 473.500 0.600 475.500 ;
    RECT 0 476.100 0.600 478.100 ;
    RECT 0 478.700 0.600 480.700 ;
    RECT 0 481.300 0.600 483.300 ;
    RECT 0 483.900 0.600 485.900 ;
    RECT 0 486.500 0.600 488.500 ;
    RECT 0 489.100 0.600 491.100 ;
    RECT 0 491.700 0.600 493.700 ;
    RECT 0 494.300 0.600 496.300 ;
    RECT 0 496.900 0.600 498.900 ;
    RECT 0 499.500 0.600 501.500 ;
    RECT 0 502.100 0.600 504.100 ;
    RECT 0 504.700 0.600 506.700 ;
    RECT 0 507.300 0.600 509.300 ;
    RECT 0 509.900 0.600 511.900 ;
    RECT 0 512.500 0.600 514.500 ;
    RECT 0 515.100 0.600 517.100 ;
    RECT 0 517.700 0.600 519.700 ;
    RECT 0 520.300 0.600 522.300 ;
    RECT 0 522.900 0.600 524.900 ;
    RECT 0 525.500 0.600 527.500 ;
    RECT 0 528.100 0.600 530.100 ;
    RECT 0 530.700 0.600 532.700 ;
    RECT 0 533.300 0.600 535.300 ;
    RECT 0 535.900 0.600 537.900 ;
    RECT 0 538.500 0.600 540.500 ;
    RECT 0 541.100 0.600 543.100 ;
    RECT 0 543.700 0.600 545.700 ;
    RECT 0 546.300 0.600 548.300 ;
    RECT 0 548.900 0.600 550.900 ;
    RECT 0 551.500 0.600 553.500 ;
    RECT 0 554.100 0.600 581.450 ;
    RECT 0 582.050 0.600 584.050 ;
    RECT 0 584.650 0.600 586.650 ;
    RECT 0 587.250 0.600 589.250 ;
    RECT 0 589.850 0.600 591.850 ;
    RECT 0 592.450 0.600 594.450 ;
    RECT 0 595.050 0.600 597.050 ;
    RECT 0 597.650 0.600 599.650 ;
    RECT 0 600.250 0.600 602.250 ;
    RECT 0 602.850 0.600 630.200 ;
    RECT 0 630.800 0.600 632.800 ;
    RECT 0 633.400 0.600 635.400 ;
    RECT 0 636.000 0.600 657.000 ;
    LAYER met4 ;
    RECT 0 0 316.800 6.500 ;
    RECT 0 650.500 316.800 657.000 ;
    RECT 0.000 6.500 5.300 650.500 ;
    RECT 7.700 6.500 10.500 650.500 ;
    RECT 12.900 6.500 15.700 650.500 ;
    RECT 18.100 6.500 20.900 650.500 ;
    RECT 23.300 6.500 26.100 650.500 ;
    RECT 28.500 6.500 31.300 650.500 ;
    RECT 33.700 6.500 36.500 650.500 ;
    RECT 38.900 6.500 41.700 650.500 ;
    RECT 44.100 6.500 46.900 650.500 ;
    RECT 49.300 6.500 52.100 650.500 ;
    RECT 54.500 6.500 57.300 650.500 ;
    RECT 59.700 6.500 62.500 650.500 ;
    RECT 64.900 6.500 67.700 650.500 ;
    RECT 70.100 6.500 72.900 650.500 ;
    RECT 75.300 6.500 78.100 650.500 ;
    RECT 80.500 6.500 83.300 650.500 ;
    RECT 85.700 6.500 88.500 650.500 ;
    RECT 90.900 6.500 93.700 650.500 ;
    RECT 96.100 6.500 98.900 650.500 ;
    RECT 101.300 6.500 104.100 650.500 ;
    RECT 106.500 6.500 109.300 650.500 ;
    RECT 111.700 6.500 114.500 650.500 ;
    RECT 116.900 6.500 119.700 650.500 ;
    RECT 122.100 6.500 124.900 650.500 ;
    RECT 127.300 6.500 130.100 650.500 ;
    RECT 132.500 6.500 135.300 650.500 ;
    RECT 137.700 6.500 140.500 650.500 ;
    RECT 142.900 6.500 145.700 650.500 ;
    RECT 148.100 6.500 150.900 650.500 ;
    RECT 153.300 6.500 156.100 650.500 ;
    RECT 158.500 6.500 161.300 650.500 ;
    RECT 163.700 6.500 166.500 650.500 ;
    RECT 168.900 6.500 171.700 650.500 ;
    RECT 174.100 6.500 176.900 650.500 ;
    RECT 179.300 6.500 182.100 650.500 ;
    RECT 184.500 6.500 187.300 650.500 ;
    RECT 189.700 6.500 192.500 650.500 ;
    RECT 194.900 6.500 197.700 650.500 ;
    RECT 200.100 6.500 202.900 650.500 ;
    RECT 205.300 6.500 208.100 650.500 ;
    RECT 210.500 6.500 213.300 650.500 ;
    RECT 215.700 6.500 218.500 650.500 ;
    RECT 220.900 6.500 223.700 650.500 ;
    RECT 226.100 6.500 228.900 650.500 ;
    RECT 231.300 6.500 234.100 650.500 ;
    RECT 236.500 6.500 239.300 650.500 ;
    RECT 241.700 6.500 244.500 650.500 ;
    RECT 246.900 6.500 249.700 650.500 ;
    RECT 252.100 6.500 254.900 650.500 ;
    RECT 257.300 6.500 260.100 650.500 ;
    RECT 262.500 6.500 265.300 650.500 ;
    RECT 267.700 6.500 270.500 650.500 ;
    RECT 272.900 6.500 275.700 650.500 ;
    RECT 278.100 6.500 280.900 650.500 ;
    RECT 283.300 6.500 286.100 650.500 ;
    RECT 288.500 6.500 291.300 650.500 ;
    RECT 293.700 6.500 296.500 650.500 ;
    RECT 298.900 6.500 301.700 650.500 ;
    RECT 304.100 6.500 306.900 650.500 ;
    RECT 309.300 6.500 316.800 650.500 ;
    LAYER OVERLAP ;
    RECT 0 0 316.800 657.000 ;
  END
END fakeram130_512x64

END LIBRARY
