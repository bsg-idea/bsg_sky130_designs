VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_64x15
  FOREIGN fakeram130_64x15 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1800.000 BY 800.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.550 0.900 18.450 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 30.150 0.900 31.050 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.750 0.900 43.650 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.350 0.900 56.250 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.950 0.900 68.850 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.550 0.900 81.450 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.150 0.900 94.050 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.750 0.900 106.650 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.350 0.900 119.250 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.950 0.900 131.850 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.550 0.900 144.450 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.150 0.900 157.050 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.750 0.900 169.650 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 181.350 0.900 182.250 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 193.950 0.900 194.850 ;
    END
  END w_mask_in[14]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 213.750 0.900 214.650 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 226.350 0.900 227.250 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 238.950 0.900 239.850 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 251.550 0.900 252.450 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 264.150 0.900 265.050 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 276.750 0.900 277.650 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 289.350 0.900 290.250 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 301.950 0.900 302.850 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 314.550 0.900 315.450 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 327.150 0.900 328.050 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 339.750 0.900 340.650 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 352.350 0.900 353.250 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 364.950 0.900 365.850 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 377.550 0.900 378.450 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 390.150 0.900 391.050 ;
    END
  END rd_out[14]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.950 0.900 410.850 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 422.550 0.900 423.450 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 435.150 0.900 436.050 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 447.750 0.900 448.650 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 460.350 0.900 461.250 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 472.950 0.900 473.850 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 485.550 0.900 486.450 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 498.150 0.900 499.050 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 510.750 0.900 511.650 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 523.350 0.900 524.250 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 535.950 0.900 536.850 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 548.550 0.900 549.450 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 561.150 0.900 562.050 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 573.750 0.900 574.650 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 586.350 0.900 587.250 ;
    END
  END wd_in[14]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 606.150 0.900 607.050 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 618.750 0.900 619.650 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 631.350 0.900 632.250 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 643.950 0.900 644.850 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 656.550 0.900 657.450 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 669.150 0.900 670.050 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 688.950 0.900 689.850 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 701.550 0.900 702.450 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 714.150 0.900 715.050 ;
    END
  END clk
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 16.200 18.000 19.800 782.000 ;
      RECT 45.000 18.000 48.600 782.000 ;
      RECT 73.800 18.000 77.400 782.000 ;
      RECT 102.600 18.000 106.200 782.000 ;
      RECT 131.400 18.000 135.000 782.000 ;
      RECT 160.200 18.000 163.800 782.000 ;
      RECT 189.000 18.000 192.600 782.000 ;
      RECT 217.800 18.000 221.400 782.000 ;
      RECT 246.600 18.000 250.200 782.000 ;
      RECT 275.400 18.000 279.000 782.000 ;
      RECT 304.200 18.000 307.800 782.000 ;
      RECT 333.000 18.000 336.600 782.000 ;
      RECT 361.800 18.000 365.400 782.000 ;
      RECT 390.600 18.000 394.200 782.000 ;
      RECT 419.400 18.000 423.000 782.000 ;
      RECT 448.200 18.000 451.800 782.000 ;
      RECT 477.000 18.000 480.600 782.000 ;
      RECT 505.800 18.000 509.400 782.000 ;
      RECT 534.600 18.000 538.200 782.000 ;
      RECT 563.400 18.000 567.000 782.000 ;
      RECT 592.200 18.000 595.800 782.000 ;
      RECT 621.000 18.000 624.600 782.000 ;
      RECT 649.800 18.000 653.400 782.000 ;
      RECT 678.600 18.000 682.200 782.000 ;
      RECT 707.400 18.000 711.000 782.000 ;
      RECT 736.200 18.000 739.800 782.000 ;
      RECT 765.000 18.000 768.600 782.000 ;
      RECT 793.800 18.000 797.400 782.000 ;
      RECT 822.600 18.000 826.200 782.000 ;
      RECT 851.400 18.000 855.000 782.000 ;
      RECT 880.200 18.000 883.800 782.000 ;
      RECT 909.000 18.000 912.600 782.000 ;
      RECT 937.800 18.000 941.400 782.000 ;
      RECT 966.600 18.000 970.200 782.000 ;
      RECT 995.400 18.000 999.000 782.000 ;
      RECT 1024.200 18.000 1027.800 782.000 ;
      RECT 1053.000 18.000 1056.600 782.000 ;
      RECT 1081.800 18.000 1085.400 782.000 ;
      RECT 1110.600 18.000 1114.200 782.000 ;
      RECT 1139.400 18.000 1143.000 782.000 ;
      RECT 1168.200 18.000 1171.800 782.000 ;
      RECT 1197.000 18.000 1200.600 782.000 ;
      RECT 1225.800 18.000 1229.400 782.000 ;
      RECT 1254.600 18.000 1258.200 782.000 ;
      RECT 1283.400 18.000 1287.000 782.000 ;
      RECT 1312.200 18.000 1315.800 782.000 ;
      RECT 1341.000 18.000 1344.600 782.000 ;
      RECT 1369.800 18.000 1373.400 782.000 ;
      RECT 1398.600 18.000 1402.200 782.000 ;
      RECT 1427.400 18.000 1431.000 782.000 ;
      RECT 1456.200 18.000 1459.800 782.000 ;
      RECT 1485.000 18.000 1488.600 782.000 ;
      RECT 1513.800 18.000 1517.400 782.000 ;
      RECT 1542.600 18.000 1546.200 782.000 ;
      RECT 1571.400 18.000 1575.000 782.000 ;
      RECT 1600.200 18.000 1603.800 782.000 ;
      RECT 1629.000 18.000 1632.600 782.000 ;
      RECT 1657.800 18.000 1661.400 782.000 ;
      RECT 1686.600 18.000 1690.200 782.000 ;
      RECT 1715.400 18.000 1719.000 782.000 ;
      RECT 1744.200 18.000 1747.800 782.000 ;
      RECT 1773.000 18.000 1776.600 782.000 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 30.600 18.000 34.200 782.000 ;
      RECT 59.400 18.000 63.000 782.000 ;
      RECT 88.200 18.000 91.800 782.000 ;
      RECT 117.000 18.000 120.600 782.000 ;
      RECT 145.800 18.000 149.400 782.000 ;
      RECT 174.600 18.000 178.200 782.000 ;
      RECT 203.400 18.000 207.000 782.000 ;
      RECT 232.200 18.000 235.800 782.000 ;
      RECT 261.000 18.000 264.600 782.000 ;
      RECT 289.800 18.000 293.400 782.000 ;
      RECT 318.600 18.000 322.200 782.000 ;
      RECT 347.400 18.000 351.000 782.000 ;
      RECT 376.200 18.000 379.800 782.000 ;
      RECT 405.000 18.000 408.600 782.000 ;
      RECT 433.800 18.000 437.400 782.000 ;
      RECT 462.600 18.000 466.200 782.000 ;
      RECT 491.400 18.000 495.000 782.000 ;
      RECT 520.200 18.000 523.800 782.000 ;
      RECT 549.000 18.000 552.600 782.000 ;
      RECT 577.800 18.000 581.400 782.000 ;
      RECT 606.600 18.000 610.200 782.000 ;
      RECT 635.400 18.000 639.000 782.000 ;
      RECT 664.200 18.000 667.800 782.000 ;
      RECT 693.000 18.000 696.600 782.000 ;
      RECT 721.800 18.000 725.400 782.000 ;
      RECT 750.600 18.000 754.200 782.000 ;
      RECT 779.400 18.000 783.000 782.000 ;
      RECT 808.200 18.000 811.800 782.000 ;
      RECT 837.000 18.000 840.600 782.000 ;
      RECT 865.800 18.000 869.400 782.000 ;
      RECT 894.600 18.000 898.200 782.000 ;
      RECT 923.400 18.000 927.000 782.000 ;
      RECT 952.200 18.000 955.800 782.000 ;
      RECT 981.000 18.000 984.600 782.000 ;
      RECT 1009.800 18.000 1013.400 782.000 ;
      RECT 1038.600 18.000 1042.200 782.000 ;
      RECT 1067.400 18.000 1071.000 782.000 ;
      RECT 1096.200 18.000 1099.800 782.000 ;
      RECT 1125.000 18.000 1128.600 782.000 ;
      RECT 1153.800 18.000 1157.400 782.000 ;
      RECT 1182.600 18.000 1186.200 782.000 ;
      RECT 1211.400 18.000 1215.000 782.000 ;
      RECT 1240.200 18.000 1243.800 782.000 ;
      RECT 1269.000 18.000 1272.600 782.000 ;
      RECT 1297.800 18.000 1301.400 782.000 ;
      RECT 1326.600 18.000 1330.200 782.000 ;
      RECT 1355.400 18.000 1359.000 782.000 ;
      RECT 1384.200 18.000 1387.800 782.000 ;
      RECT 1413.000 18.000 1416.600 782.000 ;
      RECT 1441.800 18.000 1445.400 782.000 ;
      RECT 1470.600 18.000 1474.200 782.000 ;
      RECT 1499.400 18.000 1503.000 782.000 ;
      RECT 1528.200 18.000 1531.800 782.000 ;
      RECT 1557.000 18.000 1560.600 782.000 ;
      RECT 1585.800 18.000 1589.400 782.000 ;
      RECT 1614.600 18.000 1618.200 782.000 ;
      RECT 1643.400 18.000 1647.000 782.000 ;
      RECT 1672.200 18.000 1675.800 782.000 ;
      RECT 1701.000 18.000 1704.600 782.000 ;
      RECT 1729.800 18.000 1733.400 782.000 ;
      RECT 1758.600 18.000 1762.200 782.000 ;
    END
  END vccd1
  OBS
    LAYER met1 ;
    RECT 0 0 1800.000 800.000 ;
    LAYER met2 ;
    RECT 0 0 1800.000 800.000 ;
    LAYER met3 ;
    RECT 0.900 0 1800.000 800.000 ;
    RECT 0 0.000 0.900 17.550 ;
    RECT 0 18.450 0.900 30.150 ;
    RECT 0 31.050 0.900 42.750 ;
    RECT 0 43.650 0.900 55.350 ;
    RECT 0 56.250 0.900 67.950 ;
    RECT 0 68.850 0.900 80.550 ;
    RECT 0 81.450 0.900 93.150 ;
    RECT 0 94.050 0.900 105.750 ;
    RECT 0 106.650 0.900 118.350 ;
    RECT 0 119.250 0.900 130.950 ;
    RECT 0 131.850 0.900 143.550 ;
    RECT 0 144.450 0.900 156.150 ;
    RECT 0 157.050 0.900 168.750 ;
    RECT 0 169.650 0.900 181.350 ;
    RECT 0 182.250 0.900 193.950 ;
    RECT 0 194.850 0.900 213.750 ;
    RECT 0 214.650 0.900 226.350 ;
    RECT 0 227.250 0.900 238.950 ;
    RECT 0 239.850 0.900 251.550 ;
    RECT 0 252.450 0.900 264.150 ;
    RECT 0 265.050 0.900 276.750 ;
    RECT 0 277.650 0.900 289.350 ;
    RECT 0 290.250 0.900 301.950 ;
    RECT 0 302.850 0.900 314.550 ;
    RECT 0 315.450 0.900 327.150 ;
    RECT 0 328.050 0.900 339.750 ;
    RECT 0 340.650 0.900 352.350 ;
    RECT 0 353.250 0.900 364.950 ;
    RECT 0 365.850 0.900 377.550 ;
    RECT 0 378.450 0.900 390.150 ;
    RECT 0 391.050 0.900 409.950 ;
    RECT 0 410.850 0.900 422.550 ;
    RECT 0 423.450 0.900 435.150 ;
    RECT 0 436.050 0.900 447.750 ;
    RECT 0 448.650 0.900 460.350 ;
    RECT 0 461.250 0.900 472.950 ;
    RECT 0 473.850 0.900 485.550 ;
    RECT 0 486.450 0.900 498.150 ;
    RECT 0 499.050 0.900 510.750 ;
    RECT 0 511.650 0.900 523.350 ;
    RECT 0 524.250 0.900 535.950 ;
    RECT 0 536.850 0.900 548.550 ;
    RECT 0 549.450 0.900 561.150 ;
    RECT 0 562.050 0.900 573.750 ;
    RECT 0 574.650 0.900 586.350 ;
    RECT 0 587.250 0.900 606.150 ;
    RECT 0 607.050 0.900 618.750 ;
    RECT 0 619.650 0.900 631.350 ;
    RECT 0 632.250 0.900 643.950 ;
    RECT 0 644.850 0.900 656.550 ;
    RECT 0 657.450 0.900 669.150 ;
    RECT 0 670.050 0.900 688.950 ;
    RECT 0 689.850 0.900 701.550 ;
    RECT 0 702.450 0.900 714.150 ;
    RECT 0 715.050 0.900 800.000 ;
    LAYER met4 ;
    RECT 0 0 1800.000 18.000 ;
    RECT 0 782.000 1800.000 800.000 ;
    RECT 0.000 18.000 16.200 782.000 ;
    RECT 19.800 18.000 30.600 782.000 ;
    RECT 34.200 18.000 45.000 782.000 ;
    RECT 48.600 18.000 59.400 782.000 ;
    RECT 63.000 18.000 73.800 782.000 ;
    RECT 77.400 18.000 88.200 782.000 ;
    RECT 91.800 18.000 102.600 782.000 ;
    RECT 106.200 18.000 117.000 782.000 ;
    RECT 120.600 18.000 131.400 782.000 ;
    RECT 135.000 18.000 145.800 782.000 ;
    RECT 149.400 18.000 160.200 782.000 ;
    RECT 163.800 18.000 174.600 782.000 ;
    RECT 178.200 18.000 189.000 782.000 ;
    RECT 192.600 18.000 203.400 782.000 ;
    RECT 207.000 18.000 217.800 782.000 ;
    RECT 221.400 18.000 232.200 782.000 ;
    RECT 235.800 18.000 246.600 782.000 ;
    RECT 250.200 18.000 261.000 782.000 ;
    RECT 264.600 18.000 275.400 782.000 ;
    RECT 279.000 18.000 289.800 782.000 ;
    RECT 293.400 18.000 304.200 782.000 ;
    RECT 307.800 18.000 318.600 782.000 ;
    RECT 322.200 18.000 333.000 782.000 ;
    RECT 336.600 18.000 347.400 782.000 ;
    RECT 351.000 18.000 361.800 782.000 ;
    RECT 365.400 18.000 376.200 782.000 ;
    RECT 379.800 18.000 390.600 782.000 ;
    RECT 394.200 18.000 405.000 782.000 ;
    RECT 408.600 18.000 419.400 782.000 ;
    RECT 423.000 18.000 433.800 782.000 ;
    RECT 437.400 18.000 448.200 782.000 ;
    RECT 451.800 18.000 462.600 782.000 ;
    RECT 466.200 18.000 477.000 782.000 ;
    RECT 480.600 18.000 491.400 782.000 ;
    RECT 495.000 18.000 505.800 782.000 ;
    RECT 509.400 18.000 520.200 782.000 ;
    RECT 523.800 18.000 534.600 782.000 ;
    RECT 538.200 18.000 549.000 782.000 ;
    RECT 552.600 18.000 563.400 782.000 ;
    RECT 567.000 18.000 577.800 782.000 ;
    RECT 581.400 18.000 592.200 782.000 ;
    RECT 595.800 18.000 606.600 782.000 ;
    RECT 610.200 18.000 621.000 782.000 ;
    RECT 624.600 18.000 635.400 782.000 ;
    RECT 639.000 18.000 649.800 782.000 ;
    RECT 653.400 18.000 664.200 782.000 ;
    RECT 667.800 18.000 678.600 782.000 ;
    RECT 682.200 18.000 693.000 782.000 ;
    RECT 696.600 18.000 707.400 782.000 ;
    RECT 711.000 18.000 721.800 782.000 ;
    RECT 725.400 18.000 736.200 782.000 ;
    RECT 739.800 18.000 750.600 782.000 ;
    RECT 754.200 18.000 765.000 782.000 ;
    RECT 768.600 18.000 779.400 782.000 ;
    RECT 783.000 18.000 793.800 782.000 ;
    RECT 797.400 18.000 808.200 782.000 ;
    RECT 811.800 18.000 822.600 782.000 ;
    RECT 826.200 18.000 837.000 782.000 ;
    RECT 840.600 18.000 851.400 782.000 ;
    RECT 855.000 18.000 865.800 782.000 ;
    RECT 869.400 18.000 880.200 782.000 ;
    RECT 883.800 18.000 894.600 782.000 ;
    RECT 898.200 18.000 909.000 782.000 ;
    RECT 912.600 18.000 923.400 782.000 ;
    RECT 927.000 18.000 937.800 782.000 ;
    RECT 941.400 18.000 952.200 782.000 ;
    RECT 955.800 18.000 966.600 782.000 ;
    RECT 970.200 18.000 981.000 782.000 ;
    RECT 984.600 18.000 995.400 782.000 ;
    RECT 999.000 18.000 1009.800 782.000 ;
    RECT 1013.400 18.000 1024.200 782.000 ;
    RECT 1027.800 18.000 1038.600 782.000 ;
    RECT 1042.200 18.000 1053.000 782.000 ;
    RECT 1056.600 18.000 1067.400 782.000 ;
    RECT 1071.000 18.000 1081.800 782.000 ;
    RECT 1085.400 18.000 1096.200 782.000 ;
    RECT 1099.800 18.000 1110.600 782.000 ;
    RECT 1114.200 18.000 1125.000 782.000 ;
    RECT 1128.600 18.000 1139.400 782.000 ;
    RECT 1143.000 18.000 1153.800 782.000 ;
    RECT 1157.400 18.000 1168.200 782.000 ;
    RECT 1171.800 18.000 1182.600 782.000 ;
    RECT 1186.200 18.000 1197.000 782.000 ;
    RECT 1200.600 18.000 1211.400 782.000 ;
    RECT 1215.000 18.000 1225.800 782.000 ;
    RECT 1229.400 18.000 1240.200 782.000 ;
    RECT 1243.800 18.000 1254.600 782.000 ;
    RECT 1258.200 18.000 1269.000 782.000 ;
    RECT 1272.600 18.000 1283.400 782.000 ;
    RECT 1287.000 18.000 1297.800 782.000 ;
    RECT 1301.400 18.000 1312.200 782.000 ;
    RECT 1315.800 18.000 1326.600 782.000 ;
    RECT 1330.200 18.000 1341.000 782.000 ;
    RECT 1344.600 18.000 1355.400 782.000 ;
    RECT 1359.000 18.000 1369.800 782.000 ;
    RECT 1373.400 18.000 1384.200 782.000 ;
    RECT 1387.800 18.000 1398.600 782.000 ;
    RECT 1402.200 18.000 1413.000 782.000 ;
    RECT 1416.600 18.000 1427.400 782.000 ;
    RECT 1431.000 18.000 1441.800 782.000 ;
    RECT 1445.400 18.000 1456.200 782.000 ;
    RECT 1459.800 18.000 1470.600 782.000 ;
    RECT 1474.200 18.000 1485.000 782.000 ;
    RECT 1488.600 18.000 1499.400 782.000 ;
    RECT 1503.000 18.000 1513.800 782.000 ;
    RECT 1517.400 18.000 1528.200 782.000 ;
    RECT 1531.800 18.000 1542.600 782.000 ;
    RECT 1546.200 18.000 1557.000 782.000 ;
    RECT 1560.600 18.000 1571.400 782.000 ;
    RECT 1575.000 18.000 1585.800 782.000 ;
    RECT 1589.400 18.000 1600.200 782.000 ;
    RECT 1603.800 18.000 1614.600 782.000 ;
    RECT 1618.200 18.000 1629.000 782.000 ;
    RECT 1632.600 18.000 1643.400 782.000 ;
    RECT 1647.000 18.000 1657.800 782.000 ;
    RECT 1661.400 18.000 1672.200 782.000 ;
    RECT 1675.800 18.000 1686.600 782.000 ;
    RECT 1690.200 18.000 1701.000 782.000 ;
    RECT 1704.600 18.000 1715.400 782.000 ;
    RECT 1719.000 18.000 1729.800 782.000 ;
    RECT 1733.400 18.000 1744.200 782.000 ;
    RECT 1747.800 18.000 1758.600 782.000 ;
    RECT 1762.200 18.000 1773.000 782.000 ;
    RECT 1776.600 18.000 1800.000 782.000 ;

  END
END fakeram130_64x15

END LIBRARY
