VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_64x7
  FOREIGN fakeram130_64x7 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1800.000 BY 800.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.550 0.900 18.450 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.750 0.900 43.650 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.950 0.900 68.850 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.150 0.900 94.050 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 118.350 0.900 119.250 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.550 0.900 144.450 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.750 0.900 169.650 ;
    END
  END w_mask_in[6]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 170.550 0.900 171.450 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.750 0.900 196.650 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.950 0.900 221.850 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 246.150 0.900 247.050 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 271.350 0.900 272.250 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 296.550 0.900 297.450 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 321.750 0.900 322.650 ;
    END
  END rd_out[6]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 323.550 0.900 324.450 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 348.750 0.900 349.650 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 373.950 0.900 374.850 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 399.150 0.900 400.050 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 424.350 0.900 425.250 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 449.550 0.900 450.450 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 474.750 0.900 475.650 ;
    END
  END wd_in[6]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 476.550 0.900 477.450 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 501.750 0.900 502.650 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 526.950 0.900 527.850 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 552.150 0.900 553.050 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 577.350 0.900 578.250 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 602.550 0.900 603.450 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 604.350 0.900 605.250 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 629.550 0.900 630.450 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 654.750 0.900 655.650 ;
    END
  END clk
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 16.200 18.000 19.800 782.000 ;
      RECT 45.000 18.000 48.600 782.000 ;
      RECT 73.800 18.000 77.400 782.000 ;
      RECT 102.600 18.000 106.200 782.000 ;
      RECT 131.400 18.000 135.000 782.000 ;
      RECT 160.200 18.000 163.800 782.000 ;
      RECT 189.000 18.000 192.600 782.000 ;
      RECT 217.800 18.000 221.400 782.000 ;
      RECT 246.600 18.000 250.200 782.000 ;
      RECT 275.400 18.000 279.000 782.000 ;
      RECT 304.200 18.000 307.800 782.000 ;
      RECT 333.000 18.000 336.600 782.000 ;
      RECT 361.800 18.000 365.400 782.000 ;
      RECT 390.600 18.000 394.200 782.000 ;
      RECT 419.400 18.000 423.000 782.000 ;
      RECT 448.200 18.000 451.800 782.000 ;
      RECT 477.000 18.000 480.600 782.000 ;
      RECT 505.800 18.000 509.400 782.000 ;
      RECT 534.600 18.000 538.200 782.000 ;
      RECT 563.400 18.000 567.000 782.000 ;
      RECT 592.200 18.000 595.800 782.000 ;
      RECT 621.000 18.000 624.600 782.000 ;
      RECT 649.800 18.000 653.400 782.000 ;
      RECT 678.600 18.000 682.200 782.000 ;
      RECT 707.400 18.000 711.000 782.000 ;
      RECT 736.200 18.000 739.800 782.000 ;
      RECT 765.000 18.000 768.600 782.000 ;
      RECT 793.800 18.000 797.400 782.000 ;
      RECT 822.600 18.000 826.200 782.000 ;
      RECT 851.400 18.000 855.000 782.000 ;
      RECT 880.200 18.000 883.800 782.000 ;
      RECT 909.000 18.000 912.600 782.000 ;
      RECT 937.800 18.000 941.400 782.000 ;
      RECT 966.600 18.000 970.200 782.000 ;
      RECT 995.400 18.000 999.000 782.000 ;
      RECT 1024.200 18.000 1027.800 782.000 ;
      RECT 1053.000 18.000 1056.600 782.000 ;
      RECT 1081.800 18.000 1085.400 782.000 ;
      RECT 1110.600 18.000 1114.200 782.000 ;
      RECT 1139.400 18.000 1143.000 782.000 ;
      RECT 1168.200 18.000 1171.800 782.000 ;
      RECT 1197.000 18.000 1200.600 782.000 ;
      RECT 1225.800 18.000 1229.400 782.000 ;
      RECT 1254.600 18.000 1258.200 782.000 ;
      RECT 1283.400 18.000 1287.000 782.000 ;
      RECT 1312.200 18.000 1315.800 782.000 ;
      RECT 1341.000 18.000 1344.600 782.000 ;
      RECT 1369.800 18.000 1373.400 782.000 ;
      RECT 1398.600 18.000 1402.200 782.000 ;
      RECT 1427.400 18.000 1431.000 782.000 ;
      RECT 1456.200 18.000 1459.800 782.000 ;
      RECT 1485.000 18.000 1488.600 782.000 ;
      RECT 1513.800 18.000 1517.400 782.000 ;
      RECT 1542.600 18.000 1546.200 782.000 ;
      RECT 1571.400 18.000 1575.000 782.000 ;
      RECT 1600.200 18.000 1603.800 782.000 ;
      RECT 1629.000 18.000 1632.600 782.000 ;
      RECT 1657.800 18.000 1661.400 782.000 ;
      RECT 1686.600 18.000 1690.200 782.000 ;
      RECT 1715.400 18.000 1719.000 782.000 ;
      RECT 1744.200 18.000 1747.800 782.000 ;
      RECT 1773.000 18.000 1776.600 782.000 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 30.600 18.000 34.200 782.000 ;
      RECT 59.400 18.000 63.000 782.000 ;
      RECT 88.200 18.000 91.800 782.000 ;
      RECT 117.000 18.000 120.600 782.000 ;
      RECT 145.800 18.000 149.400 782.000 ;
      RECT 174.600 18.000 178.200 782.000 ;
      RECT 203.400 18.000 207.000 782.000 ;
      RECT 232.200 18.000 235.800 782.000 ;
      RECT 261.000 18.000 264.600 782.000 ;
      RECT 289.800 18.000 293.400 782.000 ;
      RECT 318.600 18.000 322.200 782.000 ;
      RECT 347.400 18.000 351.000 782.000 ;
      RECT 376.200 18.000 379.800 782.000 ;
      RECT 405.000 18.000 408.600 782.000 ;
      RECT 433.800 18.000 437.400 782.000 ;
      RECT 462.600 18.000 466.200 782.000 ;
      RECT 491.400 18.000 495.000 782.000 ;
      RECT 520.200 18.000 523.800 782.000 ;
      RECT 549.000 18.000 552.600 782.000 ;
      RECT 577.800 18.000 581.400 782.000 ;
      RECT 606.600 18.000 610.200 782.000 ;
      RECT 635.400 18.000 639.000 782.000 ;
      RECT 664.200 18.000 667.800 782.000 ;
      RECT 693.000 18.000 696.600 782.000 ;
      RECT 721.800 18.000 725.400 782.000 ;
      RECT 750.600 18.000 754.200 782.000 ;
      RECT 779.400 18.000 783.000 782.000 ;
      RECT 808.200 18.000 811.800 782.000 ;
      RECT 837.000 18.000 840.600 782.000 ;
      RECT 865.800 18.000 869.400 782.000 ;
      RECT 894.600 18.000 898.200 782.000 ;
      RECT 923.400 18.000 927.000 782.000 ;
      RECT 952.200 18.000 955.800 782.000 ;
      RECT 981.000 18.000 984.600 782.000 ;
      RECT 1009.800 18.000 1013.400 782.000 ;
      RECT 1038.600 18.000 1042.200 782.000 ;
      RECT 1067.400 18.000 1071.000 782.000 ;
      RECT 1096.200 18.000 1099.800 782.000 ;
      RECT 1125.000 18.000 1128.600 782.000 ;
      RECT 1153.800 18.000 1157.400 782.000 ;
      RECT 1182.600 18.000 1186.200 782.000 ;
      RECT 1211.400 18.000 1215.000 782.000 ;
      RECT 1240.200 18.000 1243.800 782.000 ;
      RECT 1269.000 18.000 1272.600 782.000 ;
      RECT 1297.800 18.000 1301.400 782.000 ;
      RECT 1326.600 18.000 1330.200 782.000 ;
      RECT 1355.400 18.000 1359.000 782.000 ;
      RECT 1384.200 18.000 1387.800 782.000 ;
      RECT 1413.000 18.000 1416.600 782.000 ;
      RECT 1441.800 18.000 1445.400 782.000 ;
      RECT 1470.600 18.000 1474.200 782.000 ;
      RECT 1499.400 18.000 1503.000 782.000 ;
      RECT 1528.200 18.000 1531.800 782.000 ;
      RECT 1557.000 18.000 1560.600 782.000 ;
      RECT 1585.800 18.000 1589.400 782.000 ;
      RECT 1614.600 18.000 1618.200 782.000 ;
      RECT 1643.400 18.000 1647.000 782.000 ;
      RECT 1672.200 18.000 1675.800 782.000 ;
      RECT 1701.000 18.000 1704.600 782.000 ;
      RECT 1729.800 18.000 1733.400 782.000 ;
      RECT 1758.600 18.000 1762.200 782.000 ;
    END
  END vccd1
  OBS
    LAYER met1 ;
    RECT 0 0 1800.000 800.000 ;
    LAYER met2 ;
    RECT 0 0 1800.000 800.000 ;
    LAYER met3 ;
    RECT 0.900 0 1800.000 800.000 ;
    RECT 0 0.000 0.900 17.550 ;
    RECT 0 18.450 0.900 42.750 ;
    RECT 0 43.650 0.900 67.950 ;
    RECT 0 68.850 0.900 93.150 ;
    RECT 0 94.050 0.900 118.350 ;
    RECT 0 119.250 0.900 143.550 ;
    RECT 0 144.450 0.900 168.750 ;
    RECT 0 169.650 0.900 170.550 ;
    RECT 0 171.450 0.900 195.750 ;
    RECT 0 196.650 0.900 220.950 ;
    RECT 0 221.850 0.900 246.150 ;
    RECT 0 247.050 0.900 271.350 ;
    RECT 0 272.250 0.900 296.550 ;
    RECT 0 297.450 0.900 321.750 ;
    RECT 0 322.650 0.900 323.550 ;
    RECT 0 324.450 0.900 348.750 ;
    RECT 0 349.650 0.900 373.950 ;
    RECT 0 374.850 0.900 399.150 ;
    RECT 0 400.050 0.900 424.350 ;
    RECT 0 425.250 0.900 449.550 ;
    RECT 0 450.450 0.900 474.750 ;
    RECT 0 475.650 0.900 476.550 ;
    RECT 0 477.450 0.900 501.750 ;
    RECT 0 502.650 0.900 526.950 ;
    RECT 0 527.850 0.900 552.150 ;
    RECT 0 553.050 0.900 577.350 ;
    RECT 0 578.250 0.900 602.550 ;
    RECT 0 603.450 0.900 604.350 ;
    RECT 0 605.250 0.900 629.550 ;
    RECT 0 630.450 0.900 654.750 ;
    RECT 0 655.650 0.900 800.000 ;
    LAYER met4 ;
    RECT 0 0 1800.000 18.000 ;
    RECT 0 782.000 1800.000 800.000 ;
    RECT 0.000 18.000 16.200 782.000 ;
    RECT 19.800 18.000 30.600 782.000 ;
    RECT 34.200 18.000 45.000 782.000 ;
    RECT 48.600 18.000 59.400 782.000 ;
    RECT 63.000 18.000 73.800 782.000 ;
    RECT 77.400 18.000 88.200 782.000 ;
    RECT 91.800 18.000 102.600 782.000 ;
    RECT 106.200 18.000 117.000 782.000 ;
    RECT 120.600 18.000 131.400 782.000 ;
    RECT 135.000 18.000 145.800 782.000 ;
    RECT 149.400 18.000 160.200 782.000 ;
    RECT 163.800 18.000 174.600 782.000 ;
    RECT 178.200 18.000 189.000 782.000 ;
    RECT 192.600 18.000 203.400 782.000 ;
    RECT 207.000 18.000 217.800 782.000 ;
    RECT 221.400 18.000 232.200 782.000 ;
    RECT 235.800 18.000 246.600 782.000 ;
    RECT 250.200 18.000 261.000 782.000 ;
    RECT 264.600 18.000 275.400 782.000 ;
    RECT 279.000 18.000 289.800 782.000 ;
    RECT 293.400 18.000 304.200 782.000 ;
    RECT 307.800 18.000 318.600 782.000 ;
    RECT 322.200 18.000 333.000 782.000 ;
    RECT 336.600 18.000 347.400 782.000 ;
    RECT 351.000 18.000 361.800 782.000 ;
    RECT 365.400 18.000 376.200 782.000 ;
    RECT 379.800 18.000 390.600 782.000 ;
    RECT 394.200 18.000 405.000 782.000 ;
    RECT 408.600 18.000 419.400 782.000 ;
    RECT 423.000 18.000 433.800 782.000 ;
    RECT 437.400 18.000 448.200 782.000 ;
    RECT 451.800 18.000 462.600 782.000 ;
    RECT 466.200 18.000 477.000 782.000 ;
    RECT 480.600 18.000 491.400 782.000 ;
    RECT 495.000 18.000 505.800 782.000 ;
    RECT 509.400 18.000 520.200 782.000 ;
    RECT 523.800 18.000 534.600 782.000 ;
    RECT 538.200 18.000 549.000 782.000 ;
    RECT 552.600 18.000 563.400 782.000 ;
    RECT 567.000 18.000 577.800 782.000 ;
    RECT 581.400 18.000 592.200 782.000 ;
    RECT 595.800 18.000 606.600 782.000 ;
    RECT 610.200 18.000 621.000 782.000 ;
    RECT 624.600 18.000 635.400 782.000 ;
    RECT 639.000 18.000 649.800 782.000 ;
    RECT 653.400 18.000 664.200 782.000 ;
    RECT 667.800 18.000 678.600 782.000 ;
    RECT 682.200 18.000 693.000 782.000 ;
    RECT 696.600 18.000 707.400 782.000 ;
    RECT 711.000 18.000 721.800 782.000 ;
    RECT 725.400 18.000 736.200 782.000 ;
    RECT 739.800 18.000 750.600 782.000 ;
    RECT 754.200 18.000 765.000 782.000 ;
    RECT 768.600 18.000 779.400 782.000 ;
    RECT 783.000 18.000 793.800 782.000 ;
    RECT 797.400 18.000 808.200 782.000 ;
    RECT 811.800 18.000 822.600 782.000 ;
    RECT 826.200 18.000 837.000 782.000 ;
    RECT 840.600 18.000 851.400 782.000 ;
    RECT 855.000 18.000 865.800 782.000 ;
    RECT 869.400 18.000 880.200 782.000 ;
    RECT 883.800 18.000 894.600 782.000 ;
    RECT 898.200 18.000 909.000 782.000 ;
    RECT 912.600 18.000 923.400 782.000 ;
    RECT 927.000 18.000 937.800 782.000 ;
    RECT 941.400 18.000 952.200 782.000 ;
    RECT 955.800 18.000 966.600 782.000 ;
    RECT 970.200 18.000 981.000 782.000 ;
    RECT 984.600 18.000 995.400 782.000 ;
    RECT 999.000 18.000 1009.800 782.000 ;
    RECT 1013.400 18.000 1024.200 782.000 ;
    RECT 1027.800 18.000 1038.600 782.000 ;
    RECT 1042.200 18.000 1053.000 782.000 ;
    RECT 1056.600 18.000 1067.400 782.000 ;
    RECT 1071.000 18.000 1081.800 782.000 ;
    RECT 1085.400 18.000 1096.200 782.000 ;
    RECT 1099.800 18.000 1110.600 782.000 ;
    RECT 1114.200 18.000 1125.000 782.000 ;
    RECT 1128.600 18.000 1139.400 782.000 ;
    RECT 1143.000 18.000 1153.800 782.000 ;
    RECT 1157.400 18.000 1168.200 782.000 ;
    RECT 1171.800 18.000 1182.600 782.000 ;
    RECT 1186.200 18.000 1197.000 782.000 ;
    RECT 1200.600 18.000 1211.400 782.000 ;
    RECT 1215.000 18.000 1225.800 782.000 ;
    RECT 1229.400 18.000 1240.200 782.000 ;
    RECT 1243.800 18.000 1254.600 782.000 ;
    RECT 1258.200 18.000 1269.000 782.000 ;
    RECT 1272.600 18.000 1283.400 782.000 ;
    RECT 1287.000 18.000 1297.800 782.000 ;
    RECT 1301.400 18.000 1312.200 782.000 ;
    RECT 1315.800 18.000 1326.600 782.000 ;
    RECT 1330.200 18.000 1341.000 782.000 ;
    RECT 1344.600 18.000 1355.400 782.000 ;
    RECT 1359.000 18.000 1369.800 782.000 ;
    RECT 1373.400 18.000 1384.200 782.000 ;
    RECT 1387.800 18.000 1398.600 782.000 ;
    RECT 1402.200 18.000 1413.000 782.000 ;
    RECT 1416.600 18.000 1427.400 782.000 ;
    RECT 1431.000 18.000 1441.800 782.000 ;
    RECT 1445.400 18.000 1456.200 782.000 ;
    RECT 1459.800 18.000 1470.600 782.000 ;
    RECT 1474.200 18.000 1485.000 782.000 ;
    RECT 1488.600 18.000 1499.400 782.000 ;
    RECT 1503.000 18.000 1513.800 782.000 ;
    RECT 1517.400 18.000 1528.200 782.000 ;
    RECT 1531.800 18.000 1542.600 782.000 ;
    RECT 1546.200 18.000 1557.000 782.000 ;
    RECT 1560.600 18.000 1571.400 782.000 ;
    RECT 1575.000 18.000 1585.800 782.000 ;
    RECT 1589.400 18.000 1600.200 782.000 ;
    RECT 1603.800 18.000 1614.600 782.000 ;
    RECT 1618.200 18.000 1629.000 782.000 ;
    RECT 1632.600 18.000 1643.400 782.000 ;
    RECT 1647.000 18.000 1657.800 782.000 ;
    RECT 1661.400 18.000 1672.200 782.000 ;
    RECT 1675.800 18.000 1686.600 782.000 ;
    RECT 1690.200 18.000 1701.000 782.000 ;
    RECT 1704.600 18.000 1715.400 782.000 ;
    RECT 1719.000 18.000 1729.800 782.000 ;
    RECT 1733.400 18.000 1744.200 782.000 ;
    RECT 1747.800 18.000 1758.600 782.000 ;
    RECT 1762.200 18.000 1773.000 782.000 ;
    RECT 1776.600 18.000 1800.000 782.000 ;
  END
END fakeram130_64x7

END LIBRARY
